��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-K�趹���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�[@�qR��OMQ�bs	�Dc�c~ON<��;���Z��4d��{�
��|��Ȋ)zo1���á�rezxB���]Zb@�q�*�+
MہW��K�F��1�:�Ω�[@�qR��OMQ�bs	�Dc�c~ON<��;��� B]�pE���	x]̃Dj#^Da����M��L��O���1n��i
�z����)�,�˛D��w���旴4�����<��a��rl�ʩ{�Bfळ��)���X�$� ���jǎX������n�q��}�p� �Ñ�]�*�p�㈍x�!����Y�f��a�Z��Vb$���N[E�=����tL��	Z�G�a}CK�fC���4�O�"�F�È���_�O��<$e|��!���<< �sN۪�c�	u�~Rp�,k���%k�&ָ��sE��D�őⴔIꈸV�MT7xB2I�d�HnULkIh��:h
�[ϸ��W�A��S;CM���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�
+&�s�A�F�7���3�GXS����E@��~���($�J.���
�=W�֯��i@F�5�=h�GD�#�̔"v��ƒ)?˳R����.��ѬL�1m��+Y#_WӢۉ���2=�l����ј2��<���ħƿ�9c�I�?g�f�Jm*)�m��+���qH��ufҷGپ_s�JFAa��Bzb;ym��+r��JʅY�y��
r�(����5�����x%~Y�1�:�Ω��
�/�rD���J7"�x$�^w��ѬL�1m��+5z�P�_X�I�?g�f�L#����2=�l����ј2��<��e�IC�_�\�����@J
A��w|�<��y�~/r�I��
����&�ɬ� VU+I���ť1k�`��'p�@�I�?g�f��m�������d����1�]�Xy8��;6aJVlO/����\{F˯�+)ƍ�����b9���j}8o{:��͹ ��1�Z���=������l0��F��j�q	k���A�+3W�h+��&���$S�ݪ���[7�d|���XP����~#c!��q��f�}��Gظ0����Y%T��BPe.��xu	�>��l%i�-�M�g�����E����F��j��\w��0]%��C���M��cg�P��-��%Mό���.ӏwbk�$���7Z���(�
t�ژq���U� бb*	��|	�WI�����
L'���Xw�4��}�<�=�lx+~�v�ј�"��Z鎬�������(���`$�P.eE���lC��U�T�\ ���A����ɻ:�E�1N�By3��<�]�!���\B��V���#���L�
�����Yl���#�]�!��	Ǹ�y85��(�C)&���lC��U�T�\ �͹g}|�H���p��b��e������]�!��	Ǹ�y85���ǳ@�M�H�ɇM��lC��U�T�\ ��Tǯ�!�tӱ1R�m��+�ڔ�wV��'��s��lۛ��^�9��0�S�&�����"m�K7{�>P�2-i_���F�� �yz��$6ea�8���u�����B������k3��a������d���,�'���F�