��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-K�趹���J6�qQ��J6�qQ��J6�qQ�4��s�A�|Ԣ��g��B���������'Q�|FV;�SJ�)�Y¹w���j�Ѩ+_D)�}«^�Ԛ;Q����|�?]���p�����^��bg�Ѽ?��Q2�=W�֯�^��N�&��^˻f��	g�y���}�ZC��aNvA�;��>Oʉ�~09h�i��I�?g�fh>�F<}���U��d@��o�����\ �cG��Q�	}���bS�N1�	N�6��������t�
�-�M���w�1�l��=[���헧�d��r�6b��lY�y��
r�)�Y¹w����i��T!ix�AH�k[�^��_�)��6�$`f����om2@(?udG���s8[ZΑ� �}E+�pXTN�v��p&Hk�����qP}М��X����I�?g�fP���o7c��jp��{jϾn]�2&
8,���<0�u�P�^j��N�m��+��`�+N(�&l�v��w�#&�1�:�Ω�s8�R�	�}�����`h�ag������T��:r�g��1�:�Ω�s8�R�	�}�����`h�ag����pH��q|�C�}�M{jϾn]�w�Y��k��ı����~K�%��q��"R-��b����@k�ZV"���:��#tC������s��n�
8JA�g��%f<~�I�?g�f&:��r-,|�C�}�M{jϾn]��^���!ܞ��{H`N�jQwb�&m��+�ވΦ�'�'�0�Xb]&9%��_����(Ҝ�*���-���q.bZ�����g��:���Px?w��)�G�o���sp%r�M$�*�jQwb�&m��+������Dc�c~O�n|��sSL
��l�"�DUޑK�Ŀh���K�I�?g�f}�(g���̩r~8�ȭ��%��Gx$�r����;�(8����a�E�I�?g�f}�(g���̀:���o�2EAN5���I�?g�f}�(g���̀:���o�Yc�܎Ɉs�I�?g�f}�(g����TJ��M���%��Gx$�r����;�(8+�O!IA�⿂�Px?w���TS��g��:���Px?w��~��@�.��#=bԒB�V�x���:9�+�m��+���V�^狀=E�U�e a"����몝j@_8g!�`�(i3�a�\����9�	��%�	��El5]4 :��	��ϻIG\w:�'n�^0o_
-��[��π���{ ��*��Ũ���9����fԱ@I<��fҮ�w�Z�M�_F�k-�!�`�(i3�����5	���]���>����C��U���e�!�`�(i3��|g�Y�'���Xw�,bxqX�2�����Vc�@�Q�3������o���g��m�wR)$�Cbt�5�GR\����S���(�
t�ژq���U�UL:uۅ�յ����4��J8h���T��}����K�h90�j�b�`1���u.$���"�,�>E���TD���rs�i��s�٭��[Ø�;�x��`y�����
��I���!�qg�C�]X�.we.��xu	�`�-9v����� ����Q\�_q�b�*�K�:�"��.D!�`�(i3!�`�(i3!�`�(i3!�`�(i3$w�����=��CY�樅�ā⢔H����§�!�`�(i3!�`�(i3!�`�(i3!�`�(i3�B&�G��b<dY|a�� 	�J���"�������
��I���K���!�����E��@IE�U��`�-9v��X��)On�|�[]?=ߛ-���}�@4�tʀ4�!�`�(i3!�`�(i3!�`�(i3!�`�(i3F<����Nߕ����T��}����o�����:)!�1%�@�	^���y�"B��$I��w��,c�A�L'#���h����`y�����K*��Օ߶h��M{�jc�^�pl���G�P5Lݦ	r�!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3������c��,�.C$�#�̑����>�?���9	�ħ!�`�(i3!�`�(i3!�`�(i3!�`�(i3<�6�Q=᢯��0���0�R"6��m��3i�X��ﱍJ����=7��:�rQRт�"B��$I��w��,�$u$Yo�K3R�U���A���ܫ���׎o�|�o���/dN��<�!�`�(i3!�`�(i3!�`�(i3!�`�(i3<�6�Q=ψW��C�:����v�
� wL���jk],`nd�d�`H����I�E����F7G#+��3L��'99�q�V'�MC�p���lƀ��Ԕ�p!!v*!���OjV��!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3�沯ϕދf2^R���dv�
c�;����K��#�{0� ���M��2�����Vc}�1�9Bׄ����N�ߴ��g��m�wR)$�Cb�K��I/�˩��*����(�
t�ژq���U�JO8B�A�ɬc��WN�M�{�|L��U���B����r����!�`�(i3!�`�(i3!�`�(i3!�`�(i3I�9�T��Ҷ����S�����n�+_��l�+�+���K��I/+���G��c��Et��q���U���V9{)����S��!�oLe.��xu	���S8��y�)xʔ��O
�_�Z)|#9���s� ��<CS=e�d^�aN�By3��<�]�!���\B��V�۳a'[た��~=�L�;T?΁)���-��%M�:2QYeƈ)P<�ܓ�Ys� ��<C���D�kJN�By3��<�]�!��	Ǹ�y85�����3����VFj�F㒃��q�I�� �u4�B��ٴ���\���%�ݚ�Н�!�`�(i3!�`�(i3!�`�(i3!�`�(i3�R����ȱk�h2�<C�
�b2���HF3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3F���U	\�8U���l-;\��qq
�,0s���I<��f���nܰ��ْ5
�8��1�:�Ω��D�X�֍�G`�����m�+��
J��@�����h��>��b�b)�O��;�t�iZ]XF�IV��
�Qd��[Ya�<!�`�(i3�YV(��#�I`�p40�zɈC�4M/�S��\ʖ4��l�|���jWɆ&6�\]�x�Y�u���`=��r�)1w2xEWI�I+��<��/Ī���Z:�1�KB|1<\�$ͯ������'#u"����u��c�� ߖVz�ڵxd��QQ/�>����WI~�Ct���?�!�`�(i3"�,�>E����-��%Mό���.���|��p�G	kp^y�E����F��j��\w��0]�+���42�����Vc6�
f�L�qzʕ�a�N\�����ꢤ�Ogc����L�{"�,�>E����-��%M�rs�i�نW0��_Ma�~�Ǔ8���/��4��}�<��'��L��!�`�(i3c��Et�Y�{'%s2�ew�ۏO���qh����xc�a(􆿳�tP"7��%e��0�U+�qbp@����̰�!w���B}�w��/w~���j��3L��'9�f�NF��D�,�H���D�Ͱ�����!�`�(i3!�`�(i3!�`�(i3!�`�(i3+0$�oI�K&������f��Gm/s
9��
!�`�(i3!�`�(i3!�`�(i3!�`�(i3�� �JB��7C%��ـ��Ϝ���}b�z|w:R��̰�!�Xy|�W�E����F7G#+��3L��'9����$h������7ÎƖ�"k@:G�!D2W��!�`�(i3!�`�(i3!�`�(i3!�`�(i3M�8Z�XPt(o���xn�q�+��B	cB��!3C�4M/�S��ݡ��1��Y%T��BPe.��xu	���S8�bM� 2)G��8���/��,bxqX�2�����Vc�@�Q�3�=�<���>k� Ɓ����[;�W�@���+g^l����^����>4�q��]���>����C�x�j؀O��w���B}Yl���#�]�!����M[��Ǣ�\�2��s��+�w>���]2�y�Z鎬�������(���X{��N�a(􆿳����^��x�j؀O��{dOCe�@3Fj�a�k�]�!��	Ǹ�y85�BdC��S8a�bYSV7�pB�R�wX��^	QW�Q!r�{F��#��':E��7G#+�Ǘ0z�cUL�I��6���T�\ ��oR��m��%�э�:�rQRт�����
L'���Xw�.aX�bAKj�V��v� ����⎕�(�
t�������2%=dϖ�i�!�B����� j����nܰ��ْ5
�8��1�:�Ω��D�X�֌+.fu8�h���G!��:9�+�m��+��`�+N(�&l��5���m<d^c�y��A� �h�e�M�<��"�,�>E����-��%Mό���.Әy��j��k�lԇ�-{�!�`�(i3�1���o=�;��C��>��l%i�-���B['u!�`�(i3�E����F��j��\w��0]�7�����PM�'�ghR�P���
��3��]���c�A�L'@����g��'Uy\��x��7��S�n�(�a�x�f7﹏�T<9 =��ui|Ɏ;\w��0]ݑ���&�d�����l�x�f7﹏���
��3��]���>����CΌr���h�0!�`�(i3"�,�>E��c�r�,��Z鎬����7.~t=� ����8�%Y�����U�Q����z��l�q���U�(�6k�4d�V��*J !�`�(i3'�ʓv��ui|Ɏ;\w��0]�7�������!�qgE��Շ���z�ȃ�� ��]���>����C�(@X~�H:���������03R���7���Z鎬�������(����T��Uk���I�v��ݑ���&�d>&S�XQ� ":��v<�z�ȃ�� ��]���>����C΃�f�,�k]!�`�(i3"�,�>E���7���Z鎬�����m�讌�E�#D�����Ә�N^��#;r�����S��I�?g�f��R"N\����_�F��Ͱ�Tu��Q��}��N�p��G_/~.)��3\�R�F*}�c}��uO�b�^��\�-`����m�q�,j[�YP����Db��foW"�,�>E����-��%Mό���.�p�8��7��8�u?��I!�`�(i3c��Et�p�VU��Jp��T�����|��p�G	kp^y!�`�(i3c��Et��q���U��X�=)�H�7M���!�`�(i3��|g�Y�'���Xw�P���w�8Tʈ�Ym�ݡ��1��v�ј�"��Z鎬�������(���]�����|#9����o�t���⍽а"�,�>E����-��%Mό���.Ӂ��̰�!�Xy|�W!�`�(i3c��Et��q���U� бb*	��|	�WI!�`�(i3��|g�Y�'���Xw�������36��T�%G�D��#�]2�y�Z鎬�����	�7 �#֯���, e���TYl���#�]�!����M[��Ǣo;�Ul�|�Ƀ�?PA?e�J$b6�I��w��,c�A�L'#���h����`y���[��N��>&S�XQ� ":��v<�����
L'���Xw��ˣ�X| ���j!�`�(i3�]2�y�Z鎬����y��|�!�p�uF� y ������J�2��b���w�x���� �+��T���jB�Fg�Y씤`��p��>�B�㬊�N������>3��w��m�+��
J��@���D��L���_�L�Ȳ�V�溜��D�,�H�9� Im�����TƉ���S��������Ǜ�<�4����B�wj$g"�,�>E����\�vűhFyu���ߦ�(�M�--��wء}��9�sN�[7�d|���XP���f�ǩ�_yN���U��_�mD�ʮ�	�Qu�cx Lt�9r@�~����pL�� �[cz1�� ��X�j(�9��W0��gR� �ұ!�`�(i3!�`�(i3x�]�V��w�7qyX�񙗡��\���f���3�2�b^X�P�����"�,�>E��4];ˍH�6iQ����L?V{h�e.5��YQ�(*w��k/�z�xEQ!�`�(i3�����5	���]���>����C�C|0���!�`�(i3Y%T��BPe.��xu	�L$�����/���NM����U���e�!�`�(i3Y%T��BPe.��xu	�>��l%i�-���B['u!�`�(i3�E����F��j��\w��0]�o�t���J�g�*&��oF����-��%M�rs�i���	�>�g��U-�e�,���6+�g�G��0�ʪ%��1�����5	���]���>����C��(R\֎u�⍽аY%T��BPe.��xu	�>��l%i�-i��H�p!�`�(i3�E����F��j��\w��0]��0�&�ͭ�y{N�En�"�,�>E���TD��ό���.��D������Ҷ����SOL�V�j����(�
t�ژq���U�[��N����%O�	^���y�����
L'���Xwd�n]N�/��A����Q[R�7�%t̓�@�H�\�{\��jr�L.��7G#+��\w��0]��f�,�k]!�`�(i3"�,�>E���TD��ό���.�q�\E��0�-�`~ ��!�`�(i3c��Et�Y�{'%s^;$v�P��<�4�����6��	���`y����ꢤ�Og��P=�<�!�`�(i3�����
L'���Xw�j�7��*����V3���W��_�ړ8���/�&�<���8�t��]�'�ʪ%��1�]2�y�Z鎬����y��|�!�p�uF� y ������J�2��b���w�x���� �+��T���jB�Fg�Y씤`��p��>�B��7���
��# DY��JH3#��Aq��:9�+�m��+�<4��ˌ�ň��h��֑�/6K�R�pXTN�v��e a"����몾
�I�>y!�`�(i3,ԯ���gn��Ab�%^�;-оk�	ܷ�4D�P����JHn��z���z�O҈MA��W��g�&�0m�Q�^�y�zL͊�q���,Na�G�a���É�� �-����
c�����'��̃�����oP!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3��|R#�6�^{�����0̐p�Ѳ,�u�����e`Ez#j�?79���F�/L'��q�S<IÙ=�H%v@����fTN\;�6
�������i�±�sR�{F;�f��X��Ye�?���A���O𣧶�OZ�J�A( ����_ֲ��mŹ��C
����Ŗ6$\KʽI�����I��2m�h�_�y�H�RtV�^!�`�(i3!�`�(i3!�`�(i3!�`�(i3�q�	��cN,B�K��T�U!(��0��L�s�ޘ���m l�o��������D	��U�l>o��|�,+$\�M�ƕ�mo�0�VC ��0|]<w:����D	��U�l>o��|��س&<��3e>����C�z¡��h�'f R!�`�(i3��|g�Y�'���Xw�������펎��{5�E����F��j��\w��0]�+���42�����Vc6�
f�L�qzʕ�a�N\�����ꢤ�Ogc����L�{�����E��@IE�U����S8��y�)xʔ���6��	���`y�����
��I���!�qg�C�]X�.we.��xu	�`�-9v����� ����Q\�_q�b�*�K�:�"��.D!�`�(i3!�`�(i3!�`�(i3!�`�(i3$w�����=��CY�樅�ā⢔H����§�!�`�(i3!�`�(i3!�`�(i3!�`�(i3�B&�G��b<dY|a�� 	�J���"�������
��I���K���!�����E��@IE�U��`�-9v��X��)On�|�[]?=ߛ-���}�@4�tʀ4�!�`�(i3!�`�(i3!�`�(i3!�`�(i3F<����Nߕ����T��}����o�����:)!�1%�@�	^���y�"B��$I��w��,c�A�L'#���h����`y�����K*��Օ߶h��M{�jc�^�pl���G�P5Lݦ	r�!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3������c��,�.C$�#�̑����>�?���9	�ħ!�`�(i3!�`�(i3!�`�(i3!�`�(i3<�6�Q=᢯��0���0�R"6��m��3i�X��ﱍJ����=7��:�rQRт�"B��$I��w��,�$u$Yo�K3R�U���A���ܫ���׎o�|�o���/dN��<�!�`�(i3!�`�(i3!�`�(i3!�`�(i3<�6�Q=ψW��C�:����v�
� wL���jk],`nd�d�`H����I�E����F7G#+��3L��'99�q�V'�MC�p���lƀ��Ԕ�p!!v*!���OjV��!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3�沯ϕދf2^R���dv�
c�;����K��#�{0� ���M��2�����Vc}�1�9Bׄ����N�ߴ��g��m�wR)$�Cb�K��I/�˩��*����(�
t�ژq���U�JO8B�A�ɬc��WN�M�{�|L��U���B����r����!�`�(i3!�`�(i3!�`�(i3!�`�(i3I�9�T��Ҷ����S�����n�+_��l�+�+���K��I/+���G��c��Et��q���U���V9{)����S��!�oLe.��xu	���S8��y�)xʔ���6��	���`y�����V9{)=5.B����Y%T��BPe.��xu	�L$�����//��kOT������P��2Dg����|g�Y�'���Xw�����C���V9{)�����p������e.��xu	���S8�P?_������Cҷ��e�eO��u
�r�J�n[�n��iH�!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3{�K������K��S���6Y��y'��BSƫ6�I<��f���nܰ��ْ5
�8��1�:�Ω�s8�R�	�}����Q%b<Y�D��>3��w��m�+��
J��@���D��L���_�L�3��0I}.��dPc)y��k3��a�t�iZ]XF�IV��
�Q@���k��"�,�>E��ʆ�In��t��Q�]��-P�vȜ�[��CC��E\!��-IÙ=�H*.�PS�����k�5l�S2p�Մ�A( ����_ֲ��mŹ�[�g�DPp㧥���*�W���g�JHn��z���z�O҈��O���Ch<Q��T3�F�i�6�Ặ��Ϊ��p8/��e>����C�z¡��h�'f R!�`�(i3N�By3��<�]�!����M[��ǢR�����!�`�(i3v�ј�"��Z鎬����A��:6])2�����Vc2�����Vc߶�z7��Zr
�0�M�yObFT+V��퇇М1!�`�(i3N�By3��<�]�!��	Ǹ�y85�2�Ԡx��CyW�f�tR�wX��q�\E��0/s�1��p�E����F��j���0z�cUL��`��`�ю�������[��CC�z���a���ł�!r�dN�<@Iv��nt=:�:E��]��8|�;�Ojz���)e����|g�Y�'���Xw&�<���8�t��]�'�ʪ%��1c��Et��q���U�[��N�������lO�LYw9���TD��ό���.�:)!�1%�@�	^���y�E����F��j���0z�cUL�I��6���T�\ ��֕ߝԀ�2�����Vc2�����Vc�i�T� 둨t0����/��͈�N�˵q�׏�T#�3�["���N�DNl��Oh !6�e.��xu	�>��l%i�-��+g^l�>&S�XQ����&`���I��w��,>����C�x�j؀O��_���RQ�
Yl���#�]�!��	Ǹ�y85�2�Ԡx��CyW�f�tR�wX��^	QW�Q!r�fN�ї��q]�07G#+�Ǘ0z�cUL��`��`�ю�������[��CC�z���a�R�wX��^	QW�Q!r�{F��#��':E��7G#+�Ǘ0z�cUL�I��6���T�\ ��oR��m��%�э�:�rQRт�����
L'���Xw�.aX�bAKj�V��v� ����⎕�(�
t�������2%=dϖ�i�!�B����� j����nܰ��ْ5
�8��1�:�Ω�s8�R�	�}����pn�R��}�Dc�c~Oh���G!��:9�+�m��+�Z����y��pXTN�v��ea�;y� ����t�ؾ
�I�>y!�`�(i3;/�"���'n�^0o#�S�!fI�x���9pk�o�rM�e<�!�`�(i3;/�"���'n�^0o�0��w!�`�(i3!�`�(i3!�`�(i3!�`�(i3<�6�Q=��S&ϊD����*c�0)@�����Jm�W
i�c�r�!�`�(i3!�`�(i3!�`�(i3!�`�(i3��W�C����oP���o��e�<�Z˥�@1z�+J����+�;���;�6	(U ���*����i��>�`!�`�(i3!�`�(i3!�`�(i3!�`�(i3<�6�Q=̉���ߊΖ7:�Q�%q3 z�,�Q]�|�= � �Mt����!�`�(i3!�`�(i3!�`�(i3!�`�(i3�� л�5k
��F�2�q#O��*V<�ɔ�u�I1|�!�`�(i3!�`�(i3!�`�(i3!�`�(i3�� л��m��0m7B�Kԟ��j�釸�{�~Ǐ˨�g��!�`�(i3!�`�(i3!�`�(i3!�`�(i3�qb�S[Xx�R���-�a3�i�a�>���t��.�Չ_�9��V�9!�`�(i3!�`�(i3!�`�(i3!�`�(i3�G��
Z�g
`[~&�x$��:�e�hfH'��!���^><�B�n/a�τ,��G7��!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3eX+��f J�"e~��O��!�i�3���j�\�"����ݚ�Н�!�`�(i3!�`�(i3!�`�(i3!�`�(i3�,�-��L�}�x�6���7|)�`$��:�e�h�Ϧ^c!�6�tS���}n/a�τ,���r>�R���Xc���a��_r���⃇�����6f1�W�`t��9��V�9!�`�(i3!�`�(i3!�`�(i3!�`�(i3WPtA��ro��� zv�۲=�k2���9�����?�!�`�(i3�E����F��j��\w��0]��0�&�ͭ!�`�(i3�����5	���]���>����C���"����!�`�(i3v�ј�"��Z鎬�������!�"���O'{���O0�M��rs��扈!�`�(i3��|g�Y�'���Xw�j�7���5�%]���a(􆿳����^��p�n��!�`�(i3�]2�y�Z鎬�������(���Jם����"X��[�'i�!�q�1Ig� VU+I��vMb��s��
�C��9��ϥR�{ɟ=:�ْ5
�8��1�:�Ω�`��G���Dc�c~O1}Kط��4q������Tkd�_���n���	h��IB��XP���<����k�|�c8?-+eN7��c��;��\�vŮ�@W��C#/<���q�V�&��'�E����#3Y��P4p�ji�ШFs��X�vHޓh`����W�3�~�B�6��J���Z/���V�/��M?� g0/p�i�F�s�3�̞~%������a[�x�۶�kvɎ����9-�8���� �@��&}"	�c�o|e.��xu	���S8�
T�F�����lC��U�T�\ ���A����l��4:�CTv�ј�"��Z鎬�������(���/p���x�CyW�f�tR�wX���_F�k-�"�,�>E����-��%Mό���.��6[��u�a�*��R4��-��%Mό���.���|��pS���c,��-��%Mό���.�q�\E��0�?��Q����TD���rs�i��UQA$�U��֜��3�T�\ ����NF��]� VU+I��vMb��s��^���!ܞ��{H`Ne�7�A��Tx���� �+��T���.��Б����K��!�pXTN�v��ea�;y� ����t��X������tS���}n/a�τ,Sp�}�f60k��{U��֜��3��TG���PIÙ=�H%T��GF̧̈́��)�ܐ�ʟ�]�AZ��:I�"_��V����p{���,�#������s�0F�2�^���=���8��/��m�����W���9�uP��@)�|{eqG-}p�!�g�[��V�/��+d��;qVeE���jO$xU]c�h�����v�ј�"��Z鎬�������(���/p���x�CyW�f�tR�wX��q�\E��0� wp�R�4��-��%M�rs�i��UQA$��5�%]���a(􆿳����^��Y&X?r>*�3���f�]�!����M[��Ǣk/�z�xEQN�By3��<�]�!����M[��Ǣ&��s���qN�By3��<�]�!����M[��Ǣ���ꀍN�By3��<�]�!����M[��Ǣ@ E����Yl���#�]�!��	Ǹ�y85�;{��T�|>����n���:<��j�F����U��:9�+�m��+�ވΦ�'�'�0�Xb���{c���S��I�?g�fWg�X1����5y�$}��V�W�]�Xy8��;6aJVlO/���2�EN�@���k�� ���3�ҺIÙ=�Hr��~-���I�R���F��c��Z��}��	�d�bzP#�-������4Q��#��w21�X��|�C#/<���q��!�u�ǭ��k��?��}��7Q�� +@����������'�=�OT���0�4z�S4ٗG�D:�]��H/!�S�av>�)'l:}��Q�Ȩ�+)	Y���
Ta�~�4�k�|L����ҭٕ!! �ָ3�o�:��o�Y�#�Ez��R�>}1�l+Tf]�i�#�l�-Px���H��U��p騥]g,H�㓻lW���LWɆ&6�\]R!�!�=&0[����	�AR"WÝkˇU�Հz|��|g�Y�'���Xw�j�7����'�e���"j���b7|#9���[�л���7sI����͂��j���0z�cUL
 '&1��;�¬pX��g��U-�e�,���6+�k/�z�xEQN�By3��<�]�!����M[��Ǣ&��s���qN�By3��<�]�!����M[��Ǣ���ꀍN�By3��<�]�!����M[��Ǣ@ E����Yl���#�]�!��	Ǹ�y85�;{��T�|>����n���:<��j�F����U����ǥյ�1�:�Ω�P�p^��J���t��Dc�c~Oh���G!��:9�+�m��+F��8�ĭ��{0��d#�Dc�c~O1}Kط��4q�����]V�H7'�R�^Ƒ���E����F�'n�^0o�L��G|�7�`�4|�U�Ѯ�}t�	BH���s%
+2b�����9��]�i�xR��%�w��#�� ������!��
}��QҥF����x�Q����V�/�9
�H.�Ax.�N�K"��V�/����	c/�+��q~��z�$����Z>Ѿ��/@��_2�G@��I8����9D���o�j�0�J�vt�OF��������g2Uo�H�0�{�?Nt�!�ei�P�?��'&�s��Ia�|���+,�)��R�ᑧv0-�(4��AYpǞ��8sU��֜��3��TG���PIÙ=�H0/�+Ύ��M���R��ӟ-��[7�d|���XP�����<��no#��٠R�^Ƒ���b9�����w9�ѷ��[MD|����a��'�-��띂ii�4];ˍH�P�(e�X����4gkOq��f�}��?��[���-��%Mό���.��_F�k-�v�ј�"��Z鎬����F�71�B��O1��m<e.��xu	�>��l%i�-���6���p<��:�ҋX����>��l%i�-�[b�0<��c��Et�Y�{'%s��.|Z���I7��-5��6��	���`y����ꢤ�Og�ś� ����]�!��	Ǹ�y85��L�@��f�U����z~��6��	��k/��m#jAY4 mv���S��I�?g�f�SL�<.w[!�� Q鹯e)�Op$���{c���S��I�?g�f%��h,��;�0��'>�m�q�,�,\ަ�It�k\,آ(��7�j2����OtB!�`�(i3jݭ�F�����&]�+�Q��F���x.�Knq������E����F�Z�>)��<H�-��*����Kp&�@���k��!�`�(i3�����5	��{�OF8<z,Ҽ&��6p%�;>4�Rc��ٕ)����i3<�f�D���X���`)馢䃒����Q��K�����!�`�(i37�ܥ��2����*����i��>�`� �@"#��
}oX�4(���k�;�2M�W�Ặ��Ϊ��p8/��e>����Cx�;�x�[�л���7"�,�>E����-��%M�rs�i�jf� l�Ǜ������CyW�f�tR�wX��q�\E��0</���/�u��(�
t��Y�{'%s��.|Z���I7��-5��6��	���`y����*#�m z����Z��o�����
L'���Xw�j�7����w�K����+��dЧ^{�j����#oM|#9���Q3S�����o5��8�TD���rs�i���`�M�	=̞��>���I�Ūe�ǩ"�4s2��ԜF��g.�~R�a(􆿳�ټ*w2�56
���&~^)�E����F��j��\w��0]��b~y� �"�,�>E����-��%Mό���.�Ɏ�#���?\a��4��(�
t�ژq���U�,XG�wz#�9
4�٩�����
L'���Xw�6�:v/l����Sv�ј�"��Z鎬���������o�	�7��r�=N�By3��<�]�!����M[��Ǣ���ꀍ�����5	���]���>����C���"����Y%T��BPe.��xu	�*�QN����q�1Ig� VU+I��vMb��s����T-Q3�Y�ݬ�5����S��I�?g�f}�(g������̄'ubF��JT��k4 �	{����aҗ�(�Q�#<4^���{l�f|�ό���.���|��pe���b��o��C!T*�q���U��;���)"����}���v�ј�"��Z鎬�������Ӊ*K���j�������5	��]�!����M[��Ǣ��,m��Y%T��BPS�)37J*uc�A�L'�����=?�4���܂�^�Ҍ�"���H*Q��9�#2"Z鎬����ߘ�����B�r�������5	��]�!��	Ǹ�y85�<��GX��x�*aE���^����dxp	����<'���Xws�.*����!�`�(i3Yl���#�]�!��	Ǹ�y85�<��GX��x�*aE�fG�:�������a�=Aߕ��Z鎬����y��|�!�p��nܰ��ْ5
�8��1�:�Ω��#��,�K��ۭ�W;(q�L���N�p��G_�(����5�6ԊM$x->�A5���)5.Pf�����dJ�B�Y#�0^�� ��S�)37J*uc�A�L'��Åm�O�4���܂/븋�?��k<�v�&_K�]�!��	Ǹ�y85����!OF�u*w�A�������v���B�I��w��,c�A�L'��Åm�O�4���܂I<��f��F����U��:9�+�m��+^
s��fv����m�+��
J��@��sSL
��l�"�DUޑK	���NB����9����ۙ��\n�i�Z鎬�������(���2/
e�C�Yu*w�A�V9_=('��h�d �'���Xwd�n]N�W�R�ٶ�P �ZHA^�Xt��t-�]�Gڮ4\{Z鎬�������(���2/
e�C�Y�l�@qN=
��N�?�_u�
���)�*Y x�S$�r����;�(8S�J`�}�� VU+I��vMb��s����v����4W���f=1c� gs����'�N�Ae�#��4�gnAZ鎬�������(���2/
e�C�Yu*w�A4�3/Xδ!�`�(i3�����
L'���Xwd�n]N�7�����?�$����v�-��u��h;��!"�]��(�
t�������2�~�7���	��D܂�A�N�p��G_�(����5�6ԊM$x->��j��U�T+�S8�#��ْ5
�8��1�:�Ω��#��,�.�&�pQ0�ܩ#��E���9�ǒ,OFL}�k/�z�xEQv�ј�"��Z鎬�����X���*�Lt�2�t�����5	���]���>����C���"�����E����F��j��\w��0]����!�`�(i3c��Et�Y�{'%s2�ew����x,ɵU����I�����bn�����ឱWI��-��%Mό���.�4�3/Xδ!�`�(i3�����
L'���Xwd�n]N�?���iv���=�kJ��-4��h�]8e�0
A���J��@��sSL
��l�"�DUޑK�!EA;���q��"�$"�N�p��G_�(����5�6ԊM$x->�_��[Ǖ5.Pf�����G0P�=��2�|{	�]�!��	Ǹ�y85�� #�D�x�*aE�7�`K~���5���4	�]�!��	Ǹ�y85����!OF�l�@qN=
��N�?�_u�
���)�*Y x�S$�r����;�(8X����>x���� �+��T��#��=��va��FǼ�������@j�.(Wx*��+���)�7��r�=�o��C!T*�q���U�ЂDa��(o��0��77Ê7�E�4'���Xw�E�i�m}6	��	Mk�rN�By3��<�]�!����M[��Ǣ��,m��Y%T��BPS�)37J*uc�A�L'�����=?�4���܂�^�Ҍ�"���H*Q��9�#2"Z鎬����ߘ�����B�r�������5	��]�!��	Ǹ�y85�<��GX��x�*aE���^����dxp	����<'���Xws�.*����!�`�(i3Yl���#�]�!��	Ǹ�y85�<��GX��x�*aE�fG�:�������a�=Aߕ��Z鎬����y��|�!�p��nܰ��ْ5
�8��1�:�Ω��#��,�GkO������R���:9�+�m��+�q��.���m�����TƉ���S����j�}�I�3A�)Oq�,�S����Z�>)�ϳpJ1���مn�����-��S�<Ԣ��a�\�����Ş4=�����\{F˯�+)��KI�J�ځ�{�OF8<z,Ҽ&EfVNN�0|]<w:�x�]�V��;���Ӧ���\|Z��0[����	��cݍ�u����S�|JY%T��BPe.��xu	���S8�/ #O�)R�^Ƒ����"X��[��Q[R�7�� ߌ���E����F7G#+�Ǘ0z�cULjaGkƊ~F˯�+)�"j���b7|#9���|�au�(Z��I�V�~��TD���rs�i���`�M�	=̞��>���ԜF����am�Za(􆿳�ټ*w2�56E[��\ �����^��]���>����C����N4������[�]�!����M[��Ǣk/�z�xEQv�ј�"��Z鎬�����X���*�Lt�2�t��|g�Y�'���Xw�E�i�m}6	��	Mk�rc��Et������2�~�7���	��D܂�A�N�p��G_����(Ҝ��;�0��'>���{c���S��I�?g�fl�NAS*����*�H��m�q�,�,\ަ�Itnh'yt�;R�^Ƒ���E����F�'n�^0o����ו���E?��`�,��C����(��U��֜��3 ���3�ҺIÙ=�H�W\�o�N�Cݮ2����|�G�]R#$(��>��������	���ma�ȓl>o��|��'�njVfVi�÷�i8��4;�. � �	{��Y��
�iCN�By3��<�]�!����M[��Ǣ���ꀍc��Et��q���U��;���)"��,L�b#�ee.��xu	�`�-9v��!�`�(i3�8���&��+��(F����8���4q�\E��0le��ppȜ�]���c�A�L'��_��;w%��lC��U�T�\ ���A������U��o�TD���rs�i��~Ȃ�D�1�Z���=�"j���b7��:<��j�F����U��:9�+�m��+�Ƽ(��h�Dc�c~Oq��"�$"�N�p��G_/~.)��3\�R�F*}�c}��uO/����~r}�dPc)y��k3��a�t�iZ]XF�������̇��� +��E\!��-��7U��s7?7!* ���-N���\�v�0[����	��N�Ae�#�k/�z�xEQY%T��BPe.��xu	�>��l%i�-̇i�d�?�"�,�>E����-��%Mό���.���C7}�7��r�=��|g�Y�'���Xw�j�7����w�K��ݑ�][H5���8�R�wX�իRV�-����Cs��|g�Y�'���Xw��E�d��ЙMǿI?_�<��B��]�!����M[��Ǣշ�G!�CY%T��BPe.��xu	���S8�/ #O�)U��֜��3,0=]^	�&|#9���(@X~�H:#�<���Е�(�
t�ژq���U�[��N�霬�^����Ú���Z鎬�����	�7 �#�����g�0ˋ��I��w��,>����C��(R\֎u�3�i��7G#+��\w��0](@X~�H:�+�w>����(�
t��Y�{'%s��.|Z���ǚr��y�_��wBW��8���/�;9�".<�x���� �+��T���jB�Fg�Y씤`��p}RQaI+اy�TՄ�Dc�c~Oq��"�$"�N�p��G_/~.)��3\�R�F*}�c}��uO�Go@3w�^�������m�q�,�,\ަ�It�~V���#eI'�QFI%Ah�%4
>��`���o�:-j�!�ʺ�;[��\�v�j޽����E�4.@�A ��E+���`���o�䉌�+B����M<d_bX�>���δ V�Kx�.�H>�l땞KS�ȿ� nU���7U��s�����5jN�yYg��x�]�V��0[����	��N�Ae�#�k/�z�xEQ"�,�>E����-��%Mό���.���|��pe���b�N�By3��<�]�!����M[��Ǣ�8����"�,�>E����-��%M�rs�i���`�M�	=̞��>����� +'������݃�Q[R�7W1腰7�!�`�(i3��|g�Y�'���Xw-�}��d��2Dg��Y%T��BPe.��xu	�>��l%i�-Zs��wV�ES%Q���|g�Y�'���Xw�P���w�
�M���Y%T��BPe.��xu	�>��l%i�-I����hy�~?�2v�����
L'���Xw��E�d��ЙMǿI?2��,rL�,e.��xu	�>��l%i�-�r��f3c����L�{��|g�Y�'���Xw�j�7����'�\�n`��!��B�T�\ ��ń��,�HK���D��i��i����j��\w��0]g��	A�	N�c��|[v�ј�"��Z鎬�������(���/��A����Q[R�7�Ư�ճ�%�c��|[�����
L'���Xw�j�7��a(􆿳����^�����N4��|	�WI��(�
t�ژq���U��������:�rQRт�"B��$I��w��,>����C�Y*�Ld�!�`�(i3��(�
t�ژq���U��������B<�L�V_�"B��$I��w��,c�A�L' �oy�
!��9b�S� 7�v�ԯ��Q[R�7�D��Ø
��7��r�=�����
L'���Xw�j�7����w�K��ݑ�][H5���8�R�wX��Y�4Eb��~ߺ'^����*b.[P�{���6�l��eS:8��Ut��_k��~gj��~U��ڡP=�M:]�Idr��]��#'��;s�e�$X,��!Z㘢�TD��ό���.ӷ9lD��XH�ܲ�k?Yl���#�]�!����M[��Ǣ<���d1x�^>��y��TD���rs�i�kۜ��/�X2�B���s�_��wBW��8���/�;9�".<�x���� �+��T���jB�Fg�Y씤`��p}RQaI+k�U��OV��>3��w���(�|��s�����1�:�Ω�A��>s>;�Dc�c~O��j���