// megafunction wizard: %FIR Compiler II v11.1%
// GENERATION: XML
// fir_ramp.v

// Generated using ACDS version 11.1 173 at 2012.06.08.19:31:15

`timescale 1 ps / 1 ps
module fir_ramp (
		input  wire       clk,              //             clock_reset.clk
		input  wire       reset_n,          //       clock_reset_reset.reset_n
		input  wire       coeff_in_clk,     //       coeff_clock_reset.clk
		input  wire       coeff_in_areset,  // coeff_clock_reset_reset.reset
		input  wire [7:0] ast_sink_data,    //   avalon_streaming_sink.data
		output wire       ast_sink_ready,   //                        .ready
		input  wire       ast_sink_valid,   //                        .valid
		input  wire [1:0] ast_sink_error,   //                        .error
		output wire [9:0] ast_source_data,  // avalon_streaming_source.data
		input  wire       ast_source_ready, //                        .ready
		output wire       ast_source_valid, //                        .valid
		output wire [1:0] ast_source_error  //                        .error
	);

	fir_ramp_0002 fir_ramp_inst (
		.clk              (clk),              //             clock_reset.clk
		.reset_n          (reset_n),          //       clock_reset_reset.reset_n
		.coeff_in_clk     (coeff_in_clk),     //       coeff_clock_reset.clk
		.coeff_in_areset  (coeff_in_areset),  // coeff_clock_reset_reset.reset
		.ast_sink_data    (ast_sink_data),    //   avalon_streaming_sink.data
		.ast_sink_ready   (ast_sink_ready),   //                        .ready
		.ast_sink_valid   (ast_sink_valid),   //                        .valid
		.ast_sink_error   (ast_sink_error),   //                        .error
		.ast_source_data  (ast_source_data),  // avalon_streaming_source.data
		.ast_source_ready (ast_source_ready), //                        .ready
		.ast_source_valid (ast_source_valid), //                        .valid
		.ast_source_error (ast_source_error)  //                        .error
	);

endmodule
// Retrieval info: <?xml version="1.0"?>
//<!--
//	Generated by Altera MegaWizard Launcher Utility version 1.0
//	************************************************************
//	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//	************************************************************
//	Copyright (C) 1991-2012 Altera Corporation
//	Any megafunction design, and related net list (encrypted or decrypted),
//	support information, device programming or simulation file, and any other
//	associated documentation or information provided by Altera or a partner
//	under Altera's Megafunction Partnership Program may be used only to
//	program PLD devices (but not masked PLD devices) from Altera.  Any other
//	use of such megafunction design, net list, support information, device
//	programming or simulation file, or any other related documentation or
//	information is prohibited for any other purpose, including, but not
//	limited to modification, reverse engineering, de-compiling, or use with
//	any other silicon devices, unless such use is explicitly licensed under
//	a separate agreement with Altera or a megafunction partner.  Title to
//	the intellectual property, including patents, copyrights, trademarks,
//	trade secrets, or maskworks, embodied in any such megafunction design,
//	net list, support information, device programming or simulation file, or
//	any other related documentation or information provided by Altera or a
//	megafunction partner, remains with Altera, the megafunction partner, or
//	their respective licensors.  No other licenses, including any licenses
//	needed under any third party's intellectual property, are provided herein.
//-->
// Retrieval info: <instance entity-name="altera_fir_compiler_ii" version="11.1" >
// Retrieval info: 	<generic name="deviceFamily" value="Stratix IV" />
// Retrieval info: 	<generic name="filterType" value="Single Rate" />
// Retrieval info: 	<generic name="interpFactor" value="1" />
// Retrieval info: 	<generic name="decimFactor" value="1" />
// Retrieval info: 	<generic name="L_bandsFilter" value="All taps" />
// Retrieval info: 	<generic name="clockRate" value="100" />
// Retrieval info: 	<generic name="clockSlack" value="0" />
// Retrieval info: 	<generic name="speedGrade" value="Medium" />
// Retrieval info: 	<generic name="coeffReload" value="false" />
// Retrieval info: 	<generic name="baseAddress" value="0" />
// Retrieval info: 	<generic name="readWriteMode" value="Read/Write" />
// Retrieval info: 	<generic name="backPressure" value="false" />
// Retrieval info: 	<generic name="symmetryMode" value="Symmetrical" />
// Retrieval info: 	<generic name="delayRAMBlockThreshold" value="20" />
// Retrieval info: 	<generic name="dualMemDistRAMThreshold" value="1280" />
// Retrieval info: 	<generic name="mRAMThreshold" value="1000000" />
// Retrieval info: 	<generic name="hardMultiplierThreshold" value="-1" />
// Retrieval info: 	<generic name="inputRate" value="100" />
// Retrieval info: 	<generic name="inputChannelNum" value="1" />
// Retrieval info: 	<generic name="inputType" value="Signed Binary" />
// Retrieval info: 	<generic name="inputBitWidth" value="8" />
// Retrieval info: 	<generic name="inputFracBitWidth" value="0" />
// Retrieval info: 	<generic name="coeffSetRealValue" value="-9.78919382196E-4,0.0,-9.9805035664E-4,0.0,-0.00103783566135,0.0,-0.00110158684981,0.0,-0.00119501531175,0.0,-0.00132739522327,0.0,-0.00151371634061,0.0,-0.00177877460038,0.0,-0.00216536819859,0.0,-0.00275198370023,0.0,-0.00369487881757,0.0,-0.00534214749183,0.0,-0.00860447112625,0.0,-0.016540869863,0.0,-0.0453585747407,0.0,-0.405610412336,1.0,-0.405610412336,0.0,-0.0453585747407,0.0,-0.016540869863,0.0,-0.00860447112625,0.0,-0.00534214749183,0.0,-0.00369487881757,0.0,-0.00275198370023,0.0,-0.00216536819859,0.0,-0.00177877460038,0.0,-0.00151371634061,0.0,-0.00132739522327,0.0,-0.00119501531175,0.0,-0.00110158684981,0.0,-0.00103783566135,0.0,-9.9805035664E-4,0.0,-9.78919382196E-4" />
// Retrieval info: 	<generic name="coeffType" value="Signed Binary" />
// Retrieval info: 	<generic name="coeffBitWidth" value="12" />
// Retrieval info: 	<generic name="coeffFracBitWidth" value="12" />
// Retrieval info: 	<generic name="outType" value="Signed Binary" />
// Retrieval info: 	<generic name="outMSBRound" value="Truncation" />
// Retrieval info: 	<generic name="outMsbBitRem" value="8" />
// Retrieval info: 	<generic name="outLSBRound" value="Truncation" />
// Retrieval info: 	<generic name="outLsbBitRem" value="8" />
// Retrieval info: 	<generic name="resoureEstimation" value="1000,1200,10" />
// Retrieval info: 	<generic name="bankCount" value="1" />
// Retrieval info: 	<generic name="bankDisplay" value="0" />
// Retrieval info: </instance>
// IPFS_FILES : fir_ramp.vo
// RELATED_FILES: fir_ramp.v, altera_avalon_sc_fifo.v, auk_dspip_math_pkg_hpfir.vhd, auk_dspip_lib_pkg_hpfir.vhd, auk_dspip_avalon_streaming_controller_hpfir.vhd, auk_dspip_avalon_streaming_sink_hpfir.vhd, auk_dspip_avalon_streaming_source_hpfir.vhd, auk_dspip_roundsat_hpfir.vhd, fir_ramp_0002_rtl_wysiwyg.vhd, fir_ramp_0002_rtl.vhd, fir_ramp_0002_ast.vhd, fir_ramp_0002.vhd
