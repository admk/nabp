��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-K�趹���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω������?9|[�,HJ
Κ�P/�u�x�t���E�L#uc��WŬ�+�-ޗ(huUP���*+��`�<�R��
�n�T�+F��W��`��;�É_g�?�H�.J"����U���T���딣0&_���X0���2|	p��rw@	@us���\���Z�
ۍ���yq�`݊�|���"rG�
���}�\�.�DV	��dU�;�\��^�� ���K�}M^UQ�S��)�e
�9��Ax!P����,��*�b؏�@�~�S�`\��Yi?��n;�|-���g]����g�����fP����IL�+��ץ9�^kh�u��<��T��� �}+~�8Ó B]�pE(���B��|�o�r� �K�����)�݉|�7\F���r��RL�a)ѻtUWR����H7��7�ޑ����<��&g�7C��H��C=�)3�C����")�E�'3H��[e)�p�R\��ꫜp&C����/B!,�G�;(�B�T0�z$�}���E6sC&�gG��Hc�e$���=M��8�w'��(�D�&�〨����cZ	�M2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��~ǳ�!2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�tw:g�V|�hi��p�7��Z鎬�����R�LM��ħƿ�9c�5(��}���SaB:r���q P�^�&d�A|?_W�\I��^�َ2V�N�u�k1i�f1?�نN��_�Q�L���E�aC�h�>�N{a�9O��Yk"1/>���M[�a7Y��0�-�Dc�c~O1}Kط��4q����S��Ǵ��BR�^Ƒ���a�\����Ŵ�(??a,����\{F˯�+)�7��\����Ab�%^T_.�z0"���	��F�i�6�Ặ��Ϊ���Jjz�I�~�џ0I� X�1�x�]�V��;���Ӧ���\|Z��0[����	��N�Ae�#�뀟"�Xq<��z��}�0z�cUL�n����4���á�~O�"j���b7|#9����w,��������b3�'���Xw�j�7��;-;*�7���W��_�ړ8���/��:I�#���μeP�>���j���0z�cULjaGkƊ~F˯�+)�"j���b7|#9���{k�h�+���C�NZ鎬�������(���`$�P.eE���lC��U�T�\ ���A����{[�C`�X7G#+�Ǘ0z�cULjaGkƊ~F˯�+)�"j���b7���Øf4%6� �77Ê7�E�4'���Xw�f�VHF��>BH<M�z�]�!����M[��Ǣ�:��6�J�ҋX����>��l%i�-�|�)՜�4��{l�f|�(0̈��N���N�?�_u�-����#u��Yk"1/>���M[�a7Y��0�-�Dc�c~O������Ls�F�%ܪ���PL~΄gO�3f��*����"�Q:�{�1��q�©�����<��p����Գ+ڍ�P�西Q���Q�Q��èV!�����+�yƔ��u����L��>���	��z���AZ���$1&O�.�g3Z�j5�{�CL�x��m_�/��!N\PPE�H�b"�uQ��z/�B{�o
�s��$�Z;��|B[g�� ���S�@�
37�˱�5PM�^-q�x�l��1:�N�*�xSƏw0���D ML:�,�Xʚ@h!�`�(i3!�`�(i3fC��T����ܼY��j3��� Q�N��*lOO_Nc����L�{!�`�(i3,��O^�{	��O� m5Y��j3��� Q�N��*lOO_N�B�r��!�`�(i3,��O^�{	��O� m5Y��j3��� Q�N��*�������)�ak�m6!�`�(i3,��O^�{	��O� m5Y��j3��� Q�N��*�������,�Xʚ@h!�`�(i3,��O^�{	��O� m5'�u�uX]�Rn\�_�B�r��!�`�(i3!�`�(i3fC��T����ܼ�r����`�4,�pI�!�`�(i3!�`�(i3!�`�(i3�^,�E��HS����ݚ�Н����Y�l,r\����!�`�(i3!�`�(i3x&_FA"���@�ԗӯ��es��O!�`�(i3���gRI/,�Xʚ@h!�`�(i3!�`�(i3��q�Z�n&Y��!둿,��L�������$e����C�9Jn�+!�`�(i3!�`�(i3��x��̶�5�v����y@(8�4�!�`�(i3=���yp�.���.����!�`�(i3!�`�(i3��\��,&߰��U��f�?ǉ�=��Wʁ�Wp7�:�!�`�(i3!�`�(i3�X;p`�5�8Cl8R!�`�(i3�.��Ԕ�]��3a��!�`�(i3!�`�(i3�;�����^*�G�1�擕d�tu���ād�,������(]!�`�(i3!�`�(i3P*N�2��ҟm%��<^�d�tu���ād�,��x��B5�!�`�(i3!�`�(i3P*N�2��ҟm%��<^,\ͨ܉p������aUMf�n�Q]�����	!�`�(i3�����[h��f\k`.��J��ߟ{�����8n%d��z��BB���#��`'��e��`g��	M�D����6���0@�pgd@!�`�(i3!�`�(i3!�`�(i3xj����R��á�~O��&�C�/#�n�%G2_�ĉ�j!�`�(i3!�`�(i3-��A�sxW�O�,��L����6���ʛ�M>#�!�`�(i3!�`�(i3!�`�(i3���u�UgF˯�+)��&�C�/#�n�%,�Xʚ@h!�`�(i3!�`�(i3-��w¹��<d�,��L����6���_G��?u:�L��!�`�(i3!�`�(i3R�][[�!�`�(i3]|If">����A���I!�`�(i3!�`�(i3�O�΃S���ݚ�Н��r��SQQv�x�����D ML:�,�Xʚ@h���K�7���g��O5�!�`�(i3&�2�������ȍry��	�s�٩��$�f
%}�YmC,iguY��j3����:�"���g�Hn7�(���6����%�3��{?O��xT��ݚ�Н���#6q�Tl�������l6�	�6���I��`�i4����߈��,�ttT�ej�We��b=�Zt%��m&<g+b󆤐=�0��"��S8��#�Eע�L0�7��m�SƏw0��|3�o�%A�J�e�!�c�A�L'��䇭��L"-c����q�\E��0��A��)}��{_8�Y��=�}�Vݨf�?ǉ�=�ʸ=�Z�x�6_s/���
/���(�:�f,�c����L�{��n�T����,Wc��I�@�_&�X;p`�V�P�B�[RN�]�5'aT��3G?�d���&�a00��܀��	^��{��'��*�-�b�+�