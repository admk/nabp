��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-K�趹���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω��k�	G���%��%���UQ���?6U���T��ײ2��>���^k�/7�?1�(�c��ly[�$D֍r�	�tX�)�`���$��[dm��+@ˏ^ow�Vx���_>{������6��H4ٳ�k.w�.u���ŏ|{T%�at�3������ͧ͊�e����Us�JG�DGsc2�aB�>�;�C�l���o �����$[Z�i��%A�a��gs|�e
�9��Ax!P����9SA����q�HS�b"L]$7!����Y�f��a�Z��V2 �Q[7U�i�#!����P�>ol[�y������{S�O��<$e|����w'��1�:�Ω��k�	G���%��%���UQ���?6U���T�����\�4�sP	�b\qB�y$h��2���[emدQ�s�u�5Q�o�FS��n� F{�B*�2����_]�
K��&Tj�P�6
� �AH� K�`A���vJ�^��K+¬�I	�_�Մ�ѕ�������%"�;���
r[��<h$p<��|�	���k�8���҆�|n���:�o�E��ĕ��(�$��W��ih ��ѕ���Ϫ+2���O'{���O0�UxX�1��J'H��q�k��Y�"�+`VU���`�+N/��Fh�a~��1���VY�x��;K�:n##���Ψ�	�ǳ����c,>0�~G�6�&�^C��������{�;¬>P�2-i_��2f¬Y��RL�a)�O��u����H7�'*�O��3Q=b���{!�zg�Z�$gZߌ��h}�0�iH��L�8$�+:H뉉�V��=ƨ7K8� c��(�U����	x]̍��;��+e>�� 6V���~w���I
>��������V���8e3Z}�ax�� 5���_�xm7��(С�"pX�����U�?��+�x�8�n����Oq:m�j�{_5Jwʛ���[E�8z���U ��?��k�Jd����r�>>7�*���/���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc������2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h~09h�i�Nq�{5��]�0�lK'���Xw����Q4?���ʢ\��|�����o�3ts�JFAa��Bzb;ym��+a��ʁކ�+��T��C�NJ���1�:�Ω�*���g S��/P�p�i/-�#�����ˉ�1�:�Ω�s8�R�	�}�����ֶ�#3��������FqqDt���,��B	hI�ˋ����)��'����b]�U�IÙ=�H3���(mj7?7!* @���k��JHn��z�C�$��؍��R��j�.(Wx*�_F�k-�!�`�(i3��|g�Y�'���Xw��������lԇ�-{�N�By3��<�]�!����M[��Ǣ�8����v�ј�"��Z鎬�������(����F�dH�/�R�Ĳ4�������`y����>�w�Y�#+���G��v�ј�"��Z鎬�����	�7 �#�iK�D�b=4{W'M/��I��w��,>����C�pॻ}���E����F��j���0z�cULjaGkƊ~8����\.W^�V]��}R�wX�Ձ��̰�!w���B}�����
L'���Xw��E�d����N�DNl�@No��u��]�!����M[��Ǣ�K�&�a�*�p���@IE�U��>��l%i�-�%t̓�@��=�O��TD��ό���.Ӂ��̰�!_���RQ�
�����
L'���Xw�j�7����'�\�n`��!��B�T�\ ��Tǯ�!���\�<�dQ	���qk�ZV"���:��#tCE8�^��������3�C�p侢���I"���L~΄gO�3f��*����"�Q:�{�1k�ZV"���:��#tCE8�^��������3�C�p侢������0��7�$��Xo����HcTz�Uhw����\�v��\aьIR=���2�E~9���i�duKr�'i��g�,P�n�r��Ainv'�rC2˻����e}:���B0_�W[>���,D	�FWJ�)T�E����FT�%q���@����gG��ΉR�R��ƾ�9� �����؅�@����gG!1v!���F��6�JHn��z��ч��,1��; |�$:�c���g�,P�n��h^�+�>8
�O���|������6[7��Cҷ��ecx�S�����S8�/ #O�)U��֜��3,0=]^	�&|#9���aZ��qA�E}�%-pD�����v����<O��E�\ٿ�6�P�������M�|a)� ����35}jQ����4|�(.V���>&S�XQ���F$�T�q���U��@����gG=%� g�Vv�0q�#�7s�9���o}AM��`�������H���,>$�p�{�㘽2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc:#�c>��$O�a��Q�ڃ�)oY��o��Ca2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcZ��O��<�"��~Ǣ�)�s�ި��(R\֎u��xp�"�/�(R\֎u�
���=b�A=�n҂2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�u(����������a�=nY+�iS��g6����'J�c"0�ɠؘt�1��9�6O��B�
�ח�1F7���\�'_cG$W�1�sa��E��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����\���GW���6�o8:4�I���c�90��G��6�iI9�o«IX0F�Mf���{$�\���F�`yx�>�+X�[�G���K�k��M��K�&�a�� �^H�)P<�ܓ�Y�̢k���F�KD�Vr[/}>5��0jJ�_/�+�;�jmT�#�G�2ޟ'�5)��Z^�d��-��!��KVט$�W��7=�*��;"s�
nЯ�O��
G|1f��w���B}�����z��](g���М��^���'ƃ�3�Y�}	Vӯ)������7�Qڨn
�_�!�`�(i3�K�&�a�� �^H�״$(�>g��Ra])n#���r�����%t̓�@��0q�#��q9+t�}�;b�-�2��;�P�t�5$f��_Ub���uQL+��φ��<�6�C�9�*Q�AqeGfB��iK�D�b=\#�!V5ȑ�(R\֎u�3ח�ͣ�yaT��z��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc|9�=꨷�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc������7�,��n6�o8:4�I���c�90�Ǘa��x���8-|�D���"sS<�0�zG�������&G7�wtMMwÝ��O�~�@}?�gg�����g�Z��3��a���!@�f")u��r��'V`��b�n.����Dt��̴Hx$f��_Ub���uQL+��φ��<�6�
t����Yh��2gu�Kk���p7>Ug@����0����(R\֎u뫮�؉6�l;��ӥ�n4s1�%��W����' �Ϟ)�(����9v�j,�K?F��h� 9��n�7�Y���_j�����3p�(��i�>SOX19�-.|}�íN=]a��o���H�RtV�^���ܚ��@��f�\%���M,�ݚ�Н����F��O�VA�ڦ�c4�=~ Y���HF	��CH$�I��*�M/*�3�3CE'�ֶ>������X19�-.|}�íN=]a��o���H�RtV�^��#�a�Ą��$J�L�l:�
d������&G!�`�(i3VZ�ڋ���Y�ُC�YH�!�`�(i3�����!�`�(i3VZ�ڋ���Y�ٹ����-�!�`�(i3��Ě�����}Dq�f��k��^�1��Aݡ��d9=���u��r��;�jmT�#�(R\֎u��Gj7�uz_�mS8<�n�ݚ�Н�jCH�d*��=����h���>��[V�ݚ�Н�$f��_Ub�F�S�1 �$f��_Ub�F�S�1 �t�td���5�ŝku�������X!�`�(i3��w�`L�U5���M�����yV�a{�H������Aݡ��'����u��r��;�jmT�#�(R\֎u��Gj7�uz_�mS8<�n�ݚ�Н�jCH�d*��=����h�qB��S)��}Dq�f��	��x��ݚ�Н�jCH�d*��=����h�'i`.���}Dq�f�HN��R��bP�63Z�t�߆�p�h�M��/,�*Hx�g���-����!�`�(i3��;��L���W��7=�E㖯Hu��r��!�`�(i3��w�`L�U5���M���[ӝ��o7!�`�(i3��jVѭ@!�`�(i3���ܚ��@��f�\%����(�̚�ݚ�Н�$f��_Ub�F�S�1 �$f��_Ub�F�S�1 �t�td���5�ŝku��-��c�.!�`�(i3��w�`L�U5���M��4O���a���H������Aݡ��'����u��r��<�6�Q=ܲ�ۗ�DC�|���S9Զ�p����5��<�>VG��J�v�n�������_	
A�d�&�H�`b&�2�����d��R��Il_�Eʨ�`N/�����/�&~�xe�4�e��Vݵ,ku���>�%h��@ȥ%�+j�Tg	pT9w�[:��q��߆�p�h�M��/,�*Hx�g���-����!�`�(i3��;��L���W��7=�E㖯Hu��r��!�`�(i3��w�`L�U5���M�����yV�a{!�`�(i3��jVѭ@!�`�(i3���ܚ��@��f�\%��	�3���ݚ�Н�$f��_Ub�F�S�1 �$f��_Ub�F�S�1 �t�td���5���'��@�my$�N��ݚ�Н�����-J݉�|�T����m�ڨ�hծ?�{�XԔ�Z?�߸��S�Ȍi��<,�F!�ry�HÕ2��Ȅ&N'OVU��#6�S�T�ү",oMG~�@�S?�Pm�p�@OM.Ir�[�#��K��T��h`E�p�����E��D{%���!j������7��D��Ѓ�ݚ�Н�!�`�(i3��7I����H�^A02�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc{�-���"@�b��	��.���Y�PG�(��&Y��V�4Df���L2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��8@ʘ/k��~��/6�o8:4�I���c�90��G��6�iI9�o«IX0F�M� ��#�~C\���F�`yx�>�+X�[�G���K�k��M������V?��	�����{_8�Y��M��)=໺(ӈ���]!MuV�	�k��^�1��dc�@c�����h����^���� л����J�Q�A��p�WзBQcCs�)��S�29��|���#o�]�ʄ�;4�zu%��XW�G�<I�^$D���
�IӜ�_���ˋ�
nЯ�O�[��V���íN=]b~*��s��(R\֎u��Gj7�uz�Va�ir��[��o}@p?�]�}bu��r��t����}�����9����^�pƫ/X��-�����+Ut���T+���f��$J�L�l:�
d��n��<f���=m�n���Y'�=�P�ݚ�Н�7��u������v������f!�(�Mz�Iʜ��t���;b�-�2��;�P�t�5�� л�W�}h,?�ޫV�6�J�J��R�?`&v;�jmT�#ܲ�ۗ�DC�5��t�;��Cٯu)����bX1F#�֞q�$g�ޖ4��E��D{��-����!�`�(i3�����V?��Z���Ӳ�?��۳lU`7�X��=�HN��R��bP�63Z�t�5ߧE4��Fr��j�:����|_e=���s�p��ν(C����d�o�u�/�*c��ߡ�W&��M�φ��<�6�@a� ��fFMqlg{y����i�q,?5qM�����U��t�&P��r$ɓǃl[�Ƶ�xm��s��ݑ���&�dh����M�E�g�������(ӈ���m�r����*qA����6\�4�@�� �-j��uΜ�6Ä�Zj���
��Aݡ��d��-��!�$g�ޖ4=H����-��X� 2�!���MEʨ�`N/�<<��lp��N�DNlvr5�Dѯ���,:&�fh��[�? -��B�˒�ݚ�Н��(R\֎u�J�
�M�I� �����;b�-�2�n�l3D�.����^���'ƃ�3�Y^Md�D�fh��[�? �l�_>�O��=m�n�J3�~?��kH�RtV�^�%t̓�@���'|Fpॻ}���;�Q��:5A��p���F��O�}�	76�&�� Ӗ�t$�)�vx�qb�V�O�DܳJn����^x��v�Z��x�����)Ύ����XƤ5_��|ʡi��!�`�(i3!�`�(i3W�1�䉁�\1^O���*�f;� ��'��L��%�K��^/pӼ0��J�wzu�\G��1���~!�`�(i3��7I���;k<A���<o�;)�y�M�,!hޖ�A$�P������5d�	�+�&I(&�L��'ž1�|�'����u��r��Q� �_tt����˦G���;c���k+Q�h'�Ȝx�5W ��̫(� h�ҩ���B/�w���B}�����z��](g���М��^���'ƃ�3�Y1tSjv��H�����c�r%�o��<����M��f���'������-/a8!�`�(i3{U����Ɔ�w��kf��}Dq�f������!�`�(i3{U�����h!���|u�#�$IX�b��~$�
�:qEp�;�P�t�5fĉ>99��A0ok�����F��O�<��}�u嶫IX0F�M�c�r%����P��P���Z��W����H���,>$��:?���