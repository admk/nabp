��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-K�趹���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�s8�R�	�}����Q%b<Y�Dt-�!CB-U���T��ײ2��>���^k�/7�?1�(�c��ߘ�]��|�G��f�:��#tC��o�Rb�v �mD�?�D��L���_�L����\�Q^���������g�3��N�w	*D���y&�f��+K��[y��ڂ�1aY���~a1k��1�/lt�3� P�;��1�-���f񻲗��~o��:���F�q�\�7Y[���G:���z�t&!�ō�|'���@N1�w�0XL���. �m4�S��N������G�j����d�kⲛ���^���Gi���_,��?� �bRw�����IL�+�{Dr[��"]�Z��ހ��g�R��kF�M����h�;�~S0�>��D����r�����=�����Z�#>�MR�C�$�����{���_��qt�Y�V�� ��o�݊�V������P|�8��,\�������P����s���{Oz�IDԦ@l�3+~���Wy4p!�y'��BS�9|�x�p3�0���H��IPP������~=�L�R��|�Q�����&�q1-��h\�]΄,�H'u$�|��"t�<�֞��� ��X�pĕ�*�*-��������w�=UiwG8:b�1ҳϱ|�GJ Ւ�&�.=%)��� �i�{�Y0�6�2qq[2H�وt3����b�;`�%&��O]�lEGV`2����	��\7}�}�1JeD��0�cŮ�4s!��F؆����:�D	1d��5��Ժ����)W����T'.�>��ryІ�����mf��:6h�y�F��}���
x����g@��3ˣ��I䀜���U�R�^�WP���dIv�p��<2۱�,� �����K��mg͛�U����(1U^uh����Y�K� w�;�d���N�tכ݁=9�|Z���ߐ'�[�Z���1VU���+L��h��X�vB#|y{����P7�.yt�gU*Z9B[�^������+�ͫUz����~2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcMD��y�sY2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�#CC1X�G�ۄ��O���azhݪm����Y�{'%s#K�v]|n����f�Y!�1��8�h�� ����f�#�eM�f<�,=K�F��N��j��D���s��e�IC�_�\H�F?t�)�Y¹w�.� -��E�I�?g�f�Jm*)�m��+���qH��ufҷGپ_�	g�y�+��T��C�NJ���1�:�Ω�*���g S��/P�p����M��^�&d�A|?_W�\I��^�َ2V�N�u�k1i�f1?�نN��_�Q�L���E�aC�h�>�N{a�9Ow�Y��k��ı����~K�%��q��"R-��Sy���wɷY_GH�7����]n���E����F�Z�>)��p40�zɈ4X"��D�����ˇ ���3�ҺIÙ=�H*.�PS����vbëdP��]n���b9����r*�^�	�M�8Z�XPt.�!ŀ���g��ȝ�0����k�

gY{�o��eId�U�mu�!�`�(i3!�`�(i3!�`�(i3!�`�(i3O�^`Yk	�o%^�G@�w ��hk.�BY?�%�j���p|�4�f�5/�`g4�,�W%JHn��z���o�K�v��Ug�B�z������4-r��|ڑ�H���o���&�t.�}����F�Q���6zJ�%�撁cFẶ��Ϊ���E`�=PEoY��gνp�~Lܮ�G��C�(!���d˖*�t���Xswj!�`�(i3!�`�(i3!�`�(i3!�`�(i3<�6�Q=�Ea�7��m�]|Y2���L�3GA�\.�
��ڃ�"��E����F���8�TP����������s	IB�;�5�}�]����E����F���8�TP���{��XT}u��Q��WI~�Ct���?�!�`�(i3Y%T��BPe.��xu	�>��l%i�-��E/��FzM#��m�v�ј�"��Z鎬����A��:6])2�����Vc2�����Vc߶�z7��Zr
�0�M�yObFT+V��퇇М1!�`�(i3�����
L'���Xw�j�7���5�%]���a(􆿳����^��/$�ߺ��]��pZ�ì��|g�Y�'���Xw靤�:��D)Q7����H�N���,�t��0Q!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3�wx����ހ��g�R����!���!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3��
��`�VL�f{����߹�_|뷦R3��\���S)| ���j�����
L'���Xw�7��0�$�E�#s�@ҡ?��'o�}a�C��ݚ�Н�!�`�(i3!�`�(i3!�`�(i3!�`�(i3�uk�+ȭY&�;���dV���f����"�!T�J�g�*��/�p,��(�
t��Y�{'%s2�ew�a(􆿳��_�"ۆ�-:���h��g5]��C�
�b�s�P&"��>����!�`�(i3!�`�(i3!�`�(i3!�`�(i3&�sw'%�I���Pq/{����I����H��6Xk�scX{�X!,!�`�(i3!�`�(i3!�`�(i3!�`�(i3n���[ �p�ø��.��Ӡ�)�6��}�R�#��U_�������y�!�`�(i3��(�
t�ژq���U�Y�4Eb����"-�&<1����Y�e6�!s}6,o�}a�C�Ǐ˨�g��!�`�(i3!�`�(i3!�`�(i3!�`�(i3�5#<Z�D���� aV��w<����=��85?��k�*�1!�J�G��`�B7dԘ]2�y�Z鎬����s(Ǳ���:����v����	N.s���� �"���%a<��A��r�I�!�`�(i3!�`�(i3!�`�(i3!�`�(i3W�%kԒ�Peŋ�-�Shc,Ϸ�Kr%u���G>P���t�td���52�����Vc2�����Vcb{�o��Ш�G��g� ��^�5��^	QW�Q!r֯���,���j*(xI��w��,�$u$Yo�K�d�$;��(D��2G��
bH~��`��|��f�!�`�(i3!�`�(i3!�`�(i3!�`�(i3<�6�Q=[��l�,1B��CSkkѶ���� �TnX�g^	QW�Q!r�ԬQ�������ս��]���>����C�������PB<�L�V_��|g�Y�'���Xw�j�7���5�%]���a(􆿳����^��������P:�rQRт��|g�Y�'���Xw�����C���V9{)���ևAY%T��BPe.��xu	�L$�����//��kOT������PghR�P��|g�Y�'���Xw�j�7��a(􆿳�*Տ�*9hLx��UQ�`
Iܩ@�R���!�`�(i3!�`�(i3!�`�(i3!�`�(i3$w�����=��bv.�]�Ⳇk��8�?)���O��+Y#��6�SԎ6�r ]���f�+��T���jB�Fg�Y씤`��p�܂aQ��Dc�c~O������Ls�F�%ܪ���PL~΄gO�3f��*����"�Q:�{�1k�ZV"���:��#tC������s��Z������0��7���0@ȹ��ZBi�mR�5*%ol�ħ���$G��;�*O#���V�@M�~�������킝�wP0���O�����>�pP��^�ޑ��W��K�BE�U���q�
@�<[n^/��M`�8�s��������2�(���D<��9���W��@�A������$��Xo��/�b�P	ܷ�4D�P����Z�zL͊�q��C.W26K�~�J�� m���"u����(�ґ��:��$��Xo��� ���Lk�ȥ��}�tзq8�Ј)w�<�_N�h(����.]̌a�9D}D?�LC�Q��p��nk䅋�������z�]���,��"�Ln��S�WT�����NB����sݤd�/�Udb��X5zAo���E�{")8�*IL3#��F�7�j�2>�dט�w���-C���Cu�^���B0S�=�א=ͼ�\�vś��X&`�Kb�����=gA���_5p}w>���uS ��������s�0F�T��t��p�m~|��X�I��H�Y���4�'n�^0o��t��>e�=��?l�r�v���~��B�W��i�s��U��,��B �:��ۜ���>�8��<�V�@����gG�5�3��nS�dB�^�vtiDL��Oއ�?t},�׉é����b�����EN.'�d�6�91|�!��3��zl����b!��u���)s�?ۀB��+ H�n`5�fK�\w��0]7��"=��<D�n:3MO�`�Wi&���i%Q,$'���Xw�Y�r�7"�[�=�5x�46T`]-#��� �]_�d�٣���N N�S�.W���ۗ*�����1"e���b��d�٣���N N�S�)}���/���v䡩ثV�<�nbBI�d�٣���N N�S�)}���/����z�Ji�!�`�(i3xZ��j�
�|�x�D��	ܷ�4D�PSio���]��T�\ ��i3�|)sՀ]^U�*�!�>E-�NN&��}�WS���
�@����gG2^o�!�`^�Ad0_�S�
ut�q���U��@����gG$zv�+KX6و�cµ���U�gY�{'%s2�ew�a(􆿳���2����.���6�vhW�2�w����ƒ��2��;�d�٣��c�A�L' ��a���R�wX���7�b�������6}��=�����E����FZ鎬������_�,�� ʔ.te`�TmY>��'�Z�n�f��Z鎬������_�,�� ʔ.te`�>���Z�n�f��Z鎬�������*�n�B���_zx��.�yc�"1�#��d_7s�9���o>��l%i�-�_+H�]��3�;5 M!�`�(i3���+�J���q���U����S�B�I��
s�m�JHn��z��ч��݂W����^"4/���K䁊��l}�
�?�$ϙRl�b����aYM���Q]� _ό���.�}�
�?�#l'U:�g[-�¾L����Q]� _ό���.�}�
�?�#l'U:�g[��爤�зq8�Ј'���Xw�Y�r�7"���a�e56<^�p�y�Rv������4�]�!����w�Հ��a�e56<�:�-22�v"�,�>E���]�!���e��ƤHe�-�c���{L,8��6�P���7s�9���o>��l%i�-�_+H�]����6��8�ʪ%��1��Q]� _ό���.�}�
�?����:�`�h�� B�J���]�!����w�Հ���h��)�����X���}�CU�+vό���.� ��h���0�`xĀ����y��n`5�fK��@5���<ZJ�hEc�>*�K�ج�my�<.��2-7s�9���o>��l%i�-b!��uፀ����y����	��ܘq���U��@����gG�F�<�J��r,�U�Z鎬����s�A	��E ����7dh�?!�`�(i3�d�٣���N N�S��E ����Щ��O�*�3���g��d�٣���N N�S��E �����	(��7��E����FZ鎬�������(����F�dHP����|�J�=��?R�����!hh��C?�Q䨈��Q[R�7�_+H�]��j���H�Dȩ�v������Q]� _ό���.��7�b����pR����Υ�d[gзq8�Ј'���Xw�j�7���5�%]���a(􆿳���2����.��g#��U�,��/�T\�HP�<�d�٣��c�A�L'�����CyW�f�tR�wX��}�
�?�������P����݀�Jn,���`ό���.�}�
�?�������P�꠼*d�m��Q]� _ό���.�}�
�?���\���S)G�6�!~���Q]� _ό���.�}�
�?���\���S)CBg�Xs=���Q]� _ό���.�}�
�?�Vi� �Z$�I����Q]� _�rs�i��s�٭����D�h��T�\ ��i3�|)sՀ�i�p��+��ݫ&�b%%�E����FZ鎬�������(���Jם��C?�Q䨈��Q[R�7�����bp�Lt�2�t!�`�(i37s�9���o�jƓ�[b!��u��,�B��Z9�+	�0Dw��Ie�Pm!��p�̺���}�
�?�U�07�:�tMɶ���ns����٘�� ��`t�A~h}Nw�����������i���b�Z鎬������_�,�i�X�J�0��c�r%�[�ap�V��g���cό���.��7�b�������S��M�����ۜ��!�ό���.�}�
�?���$F@S֦O���'�DԖ��_}Ŀ~���
͵N�$Daf��pD���(�u�đ�= �U�1�&�q�Gw����\�������P����݀ ����7�o����>�/<�`A��_i}o�?A��\#���Ƹ���r����!�`�(i3!�`�(i3�"��ӌ�rg�G��0��6�a��^���H> ����)1�T��b9�� \6��.�g�G��0�T�B���э��6Bj�!�`�(i3!�`�(i3}Y;�jnc�n��`��O�W]�Jh�v��?�e0�~�zR4 :��	��g�MSG~?�d���&��D�U�2Y�s�?�6 ^��	^���y��!�=6s{\w��0]���8-|�Ds� ��<C���D�kJCw�Hm���K��I/�!��+L��o�;C2��2�w�����}o5XRpJ���QEi�:`�+P
��K��撂����~�A�qIp��K�;_j޻%202l/J@���~=�L�����3��1F#�֞qg��J�s����w�`L��9�l'N|~�.�u���r����!�`�(i3{�d"���*��c�d�hҜ����^JyR��o����>�/�<@���ل=����h��J�m�X,7<�S��#<��{��x^�2e�PB���r����!�`�(i3}Y;�jn��
��I�]�?��\f$��뺑(��U��)��S��PL��g���8��<֯���,�&ipu1n&!�`�(i3!�`�(i3!�`�(i3!�`�(i3����C=+fK/|ljq������PX6و�cµe�O��z%֯���,�L!�=�V-���+�^n=\f�5>�1x#0<-�1���%����Fg�U�D8�w��U���\���S)�;����6�����p'7TS?�A����9�O��F����{L,84a��|�&��}Dq�f���Aڬ&W럼�~=�L�����3���'����u��r��!�`�(i3�<@���ل=����h�Wsp[��X��=@'ѥ��Ra])n#���r����;�jmT�#������P�꠼*d�m1F#�֞qduP���2
�M����d9=���u��r��!�`�(i3h5���=�t���_j���Gƻ������Ɇ�5�!�`�(i3��\7�fˁ��7�|���޵.�۬gVdxQ,�K��I/��0�|�_�mS8<�n�ݚ�Н���+�t2��Lq��QF[��f�\%���}��ݚ�Н��Ra])n#]���\�x8�:
1���Ư����z��>!XM�#����+1��*Hx�g���-����!�`�(i3�D�������{
Bk	䶙%�+���q��!�`�(i3�k��^�1�K��I/z�
1���;#o�]�ʄ�
%�6W���N�Cٺ��G��Hb� h�ҩ�!�`�(i3@��( ���M/*�3��{��3���}Dq�f�՝� s�#���k$ !�`�(i3@��( ���M/*�3����3��[<�m��I�!�`�(i3�5ߧE4��!�`�(i3��Ě�����}Dq�f�
L	�\k]ǩ�/f�]�!�`�(i3�U�Z^�t� "���
w/��kOT����l��T���ӄ`^�Ad0t�;!��Q�����&G!�`�(i3�o�t����w�`L����Y� �K;��t��:!�`�(i31���~!�`�(i3@v��e��֯���,�ۿ���L��:����iW3��O�����%�������&G!�`�(i3�7����������EN.74/������.ݍ|�!�`�(i3�̢k���������P�꠼*d�m1F#�֞qduP���2
�M����'����u��r��!�`�(i3h5���=�t���_j���Gƻ������Ɇ�5�!�`�(i3��\7�fˁ��7�|���޵.�ۃVa�ir�K��I/��0�|��';��#j�ݚ�Н���+�t2��Lq��QF[��f�\%h���UZ���ݚ�Н��Ra])n#]���\�x8�:
1���Ư����z��>!XM�#����+1�;�.��1���-����!�`�(i3�D�������{
B֗M-k��%)z�
3Me!�`�(i3��jVѭ@!�`�(i3�D�������{
Bk	䶙%G�kk�!�`�(i3$f��_Ub�F�S�1 �fĉ>99��j���Gp�ݓ�W���q��n-���3��Y$�M`�K)��v�:�-22�vn��뾦�!�`�(i3,�˳�*C�����p���W�,�_sa��o���H�RtV�^����&��r��졾�g�Y�٩�����ݚ�Н���w�w:�!�`�(i3��Aڬ&W�����=��w)��
=I�^$D���������P�íN=]8k��.ͥ�H�RtV�^!�`�(i3�<@���ل=����h���}�%Dܭ��}Dq�f�՝� s�#��qX7'��֯���,�ۿ���L��:����iW3��OEʨ�`N/������&G!�`�(i3�7����������EN.74/������.ݍ|�!�`�(i3�̢k���������P�꠼*d�m�d��-��!duP���2
�M����d9=���u��r��!�`�(i3h5���=�t���_j���Gƻ��������[j!�`�(i3��\7�fˁ��7�|���޵.�ۃVa�ir�K��I/��0�|�_�mS8<�n�ݚ�Н���+�t2��Lq��QF[��f�\%�<4�sg�!�`�(i3�	��x��ݚ�Н���+�t2��Lq��QF[��f�\%�,�F��P��}Dq�f����%>�rGO�D mWN!�`�(i3�5ߧE4���ݚ�Н��ݗƩ�J��n���C!�`�(i3�U�Z^�t� "���
w/��kOT����l��T���ӄ`^�Ad0t�;!��Q�����&G!�`�(i3�o�t����w�`L����Y� �K;��t��:!�`�(i31���~!�`�(i3@v��e��֯���,�ۿ���L��:����iW3��O�����%�������&G!�`�(i3�7����������EN.74/������.ݍ|�!�`�(i3�̢k���������P�꠼*d�m1F#�֞qduP���2
�M����'����u��r��!�`�(i3h5���=�t���_j���Gƻ������Ɇ�5�!�`�(i3��\7�fˁ��7�|���޵.�ۃVa�ir�K��I/��0�|��';��#j�ݚ�Н���+�t2��Lq��QF[��f�\%h���UZ���ݚ�Н��Ra])n#]���\�x8�:
1���Ư����z��>!XM�#����+1�;�.��1���-����!�`�(i3�D�������{
B֗M-k��%)z�
3Me!�`�(i3��jVѭ@!�`�(i3�D�������{
Bk	䶙%G�kk�!�`�(i3$f��_Ub�F�S�1 �fĉ>99��j���Gp�ݓ�W���	�N�M��/�9ސt��+�t2��Lq��QF[��f�\%�,�F��P��}Dq�f��-�����5|��{+���ic)�̩ƍ2���l�?�{�X�[�g�DPp���ܐ�}��B7�Q�+ż٧���y4���;���;_��8W�w��fDiT˗=߫����L$�$G�A�FC�Р�(�V�?�d���&�����i/�/�b��+N���ˇM|�"D�K���'s� ��<C���D�kJCw�Hm���K��I/~��'vfwů��E~$�}>����ҖV��{/w1z��ӊ^�T�H�����x�����{���������EN.<��{��x� I,���Lq��QF[�b�m��He�yO�ȗ�I&�e!�`�(i3!�`�(i3�5jd�:@��( ���M/*�3��t>d��:w�٦K���r����!�`�(i3���D4FFb��8�#e��}���X��ͷ(�-�E�u�N�Lq��QF[�b�m��H3QAZ
0�1���~!�`�(i3!�`�(i3/��kOT�hҜ����^JyR���E�u�N�Lq��QF[�b�m��HԸ��S��@��( ���M/*�3�k�wS�op��
nЯ�O�!�`�(i3�%b0s�0�JcH����J�m�X,7<�S��#`H�≶�"ڊ������r����!�`�(i3}Y;�jn`���*1U�7˖�ɳ
xM�v.����U%H�(��V�j��̖UB�no�����2���:
1���ƈZeLQ��B֯���,�{W@!��e�D.7�k�#�#6��!�`�(i3!�`�(i3!�`�(i3!�`�(i3�K��I/�W[/K�W5���~=�L�����3���G�k�a�|�=�_2<:!�`�(i3!�`�(i3!�`�(i3!�`�(i3������P����/j`R�K׈
��'l/7w|]�e@��w����+�^n=\f�5>�1x#0<-�1���%�������{aO8�w��U���\���S)�;����6�����p'7TS?�A����9�O��F����{L,84a��|�&ž_�F��H�����K��I/N#~8"�Z��l[�Ƶ�1tSjv�!�`�(i3@��( ���M/*�3�c�u��nu p��@���!�`�(i3i�:`�+PN#~8"�Z�z��B��������p�:��q�՝� s�#���k$ ����l��T���ӄ��!�qgy�`��vN*���k� �ԬQ����5��t�*���k� �q� P�G��Hb� h�ҩ�!�`�(i3@��( ���M/*�3��A~����>������!�`�(i3i�:`�+PN#~8"�Z�*\�x9?&�8���&�
�:qEpm���n����7�|���޵.�ۃVa�ir�K��I/��0�|섃Va�ir�K��I/�n�{ .p�x{^4��*m!�`�(i3����&��r��졾�g��]~ڣ]�,�F��P��}Dq�f�!�`�(i3�J�g�*����3����_r��Ӝ�}Dq�f�՝� s�#���k$ !�`�(i3@��( ���M/*�3�IX�B��7��Ɇ�5�!�`�(i3T�=qއ*|X6و�cµ���(A�,"T�z�D�R!�`�(i3�5ߧE4��!�`�(i3��Ě�����}Dq�f�`���*1ʁ���MյG-0��`����>e�|����S�n�(�a����ִ��}Dq�f��-�����@:[�Xw�`v@C-�!�`�(i3,�˳�*C�����p���W�,�_sa��o���H�RtV�^����&��r��졾�g��]~ڣ]�,�F��P��}Dq�f����M$��2�w����� �.J�>��2�N�3����ۺ�u��ݚ�Н��̢k���������P�ڎC�?���v[v%���e�D.7�q���f�e�M?��y�!�`�(i3�D�������{
B��e�g��g!�%=F�=!�`�(i3:)!�1%�@�	^���yCw�Hm���B-�QŤ!�`�(i36�B��~ ��A�Y�
���3ʩ�E�1�^�
%�6W��b�3�旅Va�ir�K��I/��0�|�g�d�H�RtV�^����&��r��졾�g��]~ڣ]�,�F��P��}Dq�f����M$��2�w����� �.J�>��l8R��!�`�(i3�����!�`�(i3���g!h!�T�g�����c��۶&��L�H��>E-�N�Ӗ������%a t��e�D.7�q���f�e���v[v%������=��w)��
=a��o���H�RtV�^!�`�(i3�<@���ل=����h��{��3���}Dq�f�!�`�(i3�J�g�*����3���įէ3��}Dq�f�՝� s�#��qX7'��]�Լ�c�#o�]�ʄ����n�0R��#���n�W�G��!*���k� �ԬQ����5��t�*���k� ֯���,mk��L�������&G!�`�(i3�7����������EN.�r6���`�/{B�!�`�(i3ђw�)�WA�qIp��K/�k�2�n�)�� �g!�`�(i3�̢k�����Tյ���#���n�W�G��!*���k� �ԬQ���Kͽ<\��*���k� ֯���,mk��L�ǎ`� ܄'�!�`�(i3b��.+�s밎�+1��*Hx�g�>!XM�#�[��l�,t���H[W?ð��T�ݚ�Н���+�t2��Lq��QF[�Z9�+	�]
���7Ϝ�}Dq�f�!�`�(i3�J�g�*����3���įէ3��}Dq�f�՝� s�#W���wL�'l/7w|]�o
�Z���\(�`�����=��w)��
=
Ҥ,�㖱8�_?�b�3�怜gVdxQ,�K��I/z�
1���;����VPYu��r��!�`�(i3h5���=�t���_j���M}����BfF~X�E�ܩ<��!�`�(i3ђw�)�WA�qIp��K/�k�2�n�)�� �g!�`�(i3�̢k�����Tյ���#���n�W�G��!*���k� ]�Լ�c���J����
%�6W���N�Cٺ��#o�]�ʄ�
%�6W����!�qg�L�[\�"��-����!�`�(i3�D�������{
B��e�g��g!�%=F�=!�`�(i3���M$��2�w����� �.J�>[{�w[f!�`�(i3�	��x��ݚ�Н���+�t2��Lq��QF[�Z9�+	�Wsp[��X��=@'ѥ�!�`�(i3i�:`�+PN#~8"�Z��mU���p�8���&�
�:qEp�;�P�t�5!�`�(i3���F��O��ݚ�Н��ݗƩ��;C�T�L!�`�(i3&����aq���״$(�>g�!�`�(i3���4)c�ݘ<�̆x毘3)�:����l��T���ӄ`^�Ad0t�;!��Q�����&G!�`�(i3�o�t����w�`L�&�����~�G�kk�!�`�(i3C�4M/�Sн3y��(|v��t����~=�L�~,�H�͛�!�`�(i3��\7�f�J0i�,�L z�P��*���k� �ԬQ����5��t�1tSjv�!�`�(i3@��( ���M/*�3�c�u��nu p��@���!�`�(i3i�:`�+PN#~8"�Z��q�����8���&�Ra])n#~x]V�{���>E-�N�Ӗ������%a t���~=�L���Z<��A!>!XM�#����+1�;�.��1��B� �b��!�`�(i3�o�t����w�`L�&�����~�G�kk�!�`�(i3C�4M/�Sн3y�ܣ{�j+���X8e��e
�:qEp'{w#/ B!�`�(i3]���\�x8�Q:��?��I�^$D�����v�)y�Eh�ѮYț��N�����*���k� �ԬQ����5��t�*���k� ֯���,mk��L����ZAL�:f{�k�(F���7�|�[�A�JG��Hb� h�ҩ�!�`�(i3@��( ���M/*�3��A~����>������!�`�(i3i�:`�+PN#~8"�Z�*\�x9?&�8���&�
�:qEp���,��\���ևA�d��-��!��EJ��7o�*H��& ��0>!XM�#����+1�;�.��1�>!XM�#�[��l�,t���H[W?M?��y�!�`�(i3����&��r��졾�g��]~ڣ]�a�݌3)�!�`�(i3���M$��2�w����� �.J�>�u"����!�`�(i3�߆�p�h�M���yt7�o�*H��& ��0>!XM�#����+1��*Hx�g���S��>!XM�#�[��l�,t���H[W?�>Jj:&ֲ!�`�(i3�A!���iW3��O�����%����:�������7�|���޵.��g�d�H�RtV�^!�`�(i3�<@���ل=����h�s��m�Eq�e>%����!�`�(i3i�:`�+PN#~8"�Z�*\�x9?&�8���&�
�:qEp��`�ҪJ�F�z�>�/�a�'�Zy.
�@�����K��I/z�
1���;}2��L�)6g����O�Q:��?��I�^$D���������P�꠼*d�m����xQ�1tSjv�!�`�(i3�o�t����w�`L�&�����~��%���!�`�(i3!�`�(i3!�`�(i3�ǐU
���F�}қ~�!�`�(i3T�=qއ*|X6و�cµ���(A�,"T�z�D�R!�`�(i36�B��~ ��A�Y�
���3ʩ�V$=�b�������PLm�<o�̱�	P �a��e�D.7�q���f�e���v[v%������=��w)��
=I/��\]� h�ҩ�!�`�(i3@��( ���M/*�3�c�u��nu p��@���!�`�(i3C�4M/�Sн3y�ܣ{�j+�f����It�!�`�(i3��jVѭ@!�`�(i3�D�������{
B��e�g��g!�%=F�=!�`�(i3���M$��2�w����� �.J�>��l8R��!�`�(i3HN��R��bP�63Z�t���%>�rG�@�	������6��Ͳ�h"QU&U�)j�S���vo� ��M�#'�^����VA�ڦ�c4��Aڬ&W럼�~=�L�����3���'����u��r��!�`�(i3�<@���ل=����h����3��[<�m��I�!�`�(i3�J�g�*����3��?�4V�I~$�}>����=@'ѥ��Ra])n#���r����;�jmT�#������P�꠼*d�m�d��-��!duP���2
�M����d��-��!duP���2��'��a��o���H�RtV�^!�`�(i3�<@���ل=����h��{��3���}Dq�f�!�`�(i3�J�g�*����3���įէ3��}Dq�f�՝� s�#��!7�������+1�;�.��1�>!XM�#�=5.B��������xQ�1tSjv�!�`�(i3�o�t����w�`L�&�����~�G�kk�!�`�(i3ђw�)�WA�qIp��K/�k�2�]�u��y!�`�(i3��w�w:�!�`�(i3����&��r��졾�g��]~ڣ]���}��ݚ�Н��q�9�ͭ�Ƀ�?PA�g�+C��sJ�A7���ݚ�Н�fĉ>99��A0ok��
�:qEp�;�P�t�5��6��+m��o����?c$��!�`�(i3�B�+2��;�P����|e"�H�����K��I/N#~8"�Z��l[�Ƶ�1tSjv�!�`�(i3@��( ���M/*�3�c�u��nu p��@���!�`�(i3i�:`�+PN#~8"�Z�z��B��������p�:��q�՝� s�#���k$ ����l��T���ӄ��!�qgy�`��vN*���k� �ԬQ����5��t�*���k� �q� P�G��Hb� h�ҩ�!�`�(i3@��( ���M/*�3��A~����>������!�`�(i3i�:`�+PN#~8"�Z�*\�x9?&�8���&�
�:qEpm���n����7�|���޵.�ۃVa�ir�K��I/��0�|섃Va�ir�K��I/�n�{ .p�x{^4��*m!�`�(i3����&��r��졾�g��]~ڣ]�,�F��P��}Dq�f�!�`�(i3�J�g�*����3����_r��Ӝ�}Dq�f�՝� s�#���k$ !�`�(i3@��( ���M/*�3�IX�B��7��Ɇ�5�!�`�(i3T�=qއ*|X6و�cµ���(A�,"T�z�D�R!�`�(i3�5ߧE4��!�`�(i3��Ě�����}Dq�f����'��@�my$�N���ڦ`�C>fĉ>99��|��3�W?�;�끶���A��
���||�T^�����¦���7�`K~�� ӥ�hsy[6�o8:4�I���c�90Mj�dL�d�G}%����3fq�M�/�e���ɯ;xjzӝ���w3��׍�&�U��f�!�`�(i3��Bf����{_8�Y��=�}�Vݨ��}Dq�f���꼲x���՜�%P�&�t.�}�;b�-�2�tiND�S���/9�=eSe.��a��o��ѵ��.�~<�Ɵe�*|�÷�Wе !�`�(i3�'ž1�|�XƤ5_�a��o���H�RtV�^uD�*'�'DV���b�z'hۉ)��d�7�q�՝� s�#���k$ �H����6�_ܸy^��ۥ`�M?��y�!�`�(i3���l%�C3�'�c����D����:�T�p��;�{������l��ͱz�4��9���u����:�T�8�fk!�`�(i3+��/�6�.e:q|+���aY���W՝� s�#���k$ ~�vE�sy����D�� �v��}Dq�f���Ě�����}Dq�f�CQ3�u��H��̣���*ȑs��-����!�`�(i3/w1z��ӊ��<���#�b��~$�!�`�(i3�����!�`�(i3�����ya�E�Rq���my$�N��o�/���;!�`�(i3$f��_Ub�F�S�1 ����aR�!�`�(i3��Ě�����}Dq�f���Ě�����}Dq�f��5ߧE4��HN��R���IX0F�M�� �R�P9d^\'@��F�z�>�/~�[��+��/�6�.���:�s������,�ǰ����ԫ�`RO���֑5�i�Q�e	�D�6I^���9������y�l��φ��<�6�@a� ����C�'�ąd�G}%����3f��gmJ/���'ž1�|��P�:k& ��-�����D�������f�\%���}�����@|��璓�c�������t �[l;M?��yЩ���&��K�~��%5������{
BF����c����F��O�\E�W��4b����A���K�h�[e4��f"�	�D�6I^ܡ�C�\�8�o�fy�U��)���Y;e�iK-pm!9�>��n4s1�U��B��-��^�uJ#��r$ɓǉ�.y�U=������&G�7����׌�yt��\�g2�I�7�js�і��D�̢k���"��w6�0��ɗ��zi#Y)M���Fe��-�����D�����.��NM$x�p��^@ ��\�&ɖ��_j���?\�z?Xk��;�P�t�5�׹���& d��ܡ�C�\�8o�@' zSL&������_�KA]H {��u��]'\gWg��	�Z�kfcj��r���iI9�o��5�:��\���F�`y������T�8k��.ͥ�H�RtV�^�J�g�*-c[�����u"���ܹ߆�p�hؽ!�M��9�a>*<UB3 �~k�%�������&Gђw�)�WA�qIp��K�Z�-Q�L5�Ƀ�?PAA�Pz>ShR}�	76�&�� Ӗ�t$�)�vx�(����i�2�w����
��I#��2�w��������X::8���SY�N��&Y��V��ht��R����A$�P��O�@יߌ��omq�:Fa�7����os�鮊��h��<���"sS<GYqcHTX�';��#jׇӭ��3�;5 M!�`�(i3�q9+t�}�����������=�t��ܜ�[�)P<�ܓ�Y�7���������Us��O*m]/��kOTs� ��<C���f�r�w ����7����|e"������P�8�>�}��q9+t�}����@|����^a�nu4Bޗ��jw�	��ׇӭ��3�;5 M!�`�(i3'�^���������������=�t��ܜ�[���2�N�3���!�qg+�dr�����o�t��{��b�b�*q����`U�m���d�����W�^	QW�Q!r�TmY>��'(|v��t�'���>;#��򴶽!����C=+f3�{~��uz��B������ևA�E�i�m}6O�D mWN��ܐ�}Ĳ�y��iE��˼S����`����#QU�0��IuA]C��JJ�C�G����]'\gWg��	�Z�kfc�_	�Ƽ��S�J\7rc^Y�G?������t�r�"���\���F�`yx�>�+X�M?��yЮ_��>νr��U�,��/3�|* ���dN�<@Iv��nt=:�$r�t�}ik+Q�h'�Ȝx�5W ��̫(� h�ҩ��;�%�R���I�zӯ�_�mS8<�n�ݚ�Н�������P����A@z��B�������S����+Ut������F��O�}�	76�&�� Ӗ�t$�)�vx1x#0<-�1�}��u@:q��_N��K��I/H^��Ƨ�0������P�꠼*d�muK��zk��^́|�A0��d`������U��
t��I�؉P}�#�����K��I/G�?-�D,��	J��!H�N(�gOx���C+�!���;����K�I��+0◤�T�_��>���<�����%8����`���UKr��c�� �n}沁2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 �@���rah�v�G�=�4��:"��A���r!B����n��4�A��mn�ܠh��A�E'��BH��d��^ &��� tY�g�8�Ϯ�~38C��ەaY|`Ŷ�ե��{���L�S#���J����La�Nc"Mh��S(���c�1�f2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����x�D���������	��6zJ�(�sM$�'[��7%^G3�ai����BY�B��TC,o��.}�՜�w9���י!*N��nk��~��/6�o8:4�I���c�90��G��6�iI9�o«IX0F�M�@�A�KR2G�,��R(bs��2[�a��o�����]�KS�)Յ�N��I~F2�~)P<�ܓ�Y����������**,n��;c���k+Q�h'�Ȝx�5W ��̫(� h�ҩ�#l'U:�g[�x�~�߹#l'U:�g[첖�7�H)-|��Y��VF�˷��'�����j��c�Q�;�jmT�#](ùy�;��S�6����ˇ�J��&x� h�ҩ΄���������**,nI��
s�m�����M�
�:qEp'{w#/ B!�`�(i3I��
s�m�^օ?D^�։��%>�rGO�D mWNHN��R��bP�63Z�t�5ߧE4��Fr��j���_J��`CE՟y]5&��(��u������y��.T�Vَφ��<�6�@a� ��fFMqlg���+�^n=\f�5>���!$�(L�-"�(�ES�a��A(�c���_G��Hb�S���⫦��=7�ŏ�ʳ�(�)P<�ܓ�Y`��v
K<߲�1V�L�q9+t�}֖�߾�0�ʂ�j�Ï��	�l�lM�3 ԫ[=�.n��c,;?5�R�<<�U#o�]�ʄ��.�L�oDy���Բ�5��X1tSjv�`��v
K<�Y�|�8�q9+t�}�ݚ�Н��1!�J�G�W�^�|��/��kOT;�jmT�#](ùy�;U���ڑ�H�RtV�^n62�}�����\�Xn��뾦�!�`�(i3���F��O��ݚ�Н��%�r���ڣ�	���	ܷ�4D�P���?L�ܚ�-����!�`�(i3r��c��Z�_v(���?D�8��fĉ>99��A0ok��HN��R��bP�63Z�t���F��O�i ���=��IX0F�M�����y��ĥ�A�t����M~V��	��y ��f"�D�����|ag��6���r�����k6m.J�@�k�pqi���+��X0���_r�e~5�O�%E#P�����y�`��w9��x�i8B23`���x{6��H��q4\%��t�O��-q#λ��$��]�N��+8H{^��/!Z��E��3?�d���&�Z�7� �o�x���!�`�(i3!�`�(i3!�`�(i3��+öz��X�bJ�u8z�����X���Kp��^�#λ��$��]�N��+
‮H){�x_�o����!�5��N?g���Ο��ٴܻ�@`u:j1�e�ǦU��֜��3�9�Ek9ԔY�|�8KZ	��\#�!�`�(i3&b����H#λ��$��]�N��+"j���b7���Øf�8��N�,Ou�X#*ݔL���}ؗO=�W��H�Ů�n/��Ƀ�?PA�9*�Mmh�9�sm���}0[�d{��>[��s�A>��R{	�rO�0|�d��_��=�3��3R�>Tr*؄�N��y�@���i�{d��L��>P�֌d {�>����5i�i�ѓ;% ���W���f� �� 2����Ă�78�T��8x����c����*��gg���yM�����)��}0[�fA~,���f+��hg�>ӾӉV�ͥ$�za��B�&���oH^���rU��c,g�vG[o⷟L*��v���bQ�*�8��	�D�6I^(�"x6�if*� ��o%ˡ�؞h���m���d����Ў��:
1����r��x�~̖UB�no�^�q���j�p�U�07�:�;#�]�g����n4s1�U��B��-��& d��]�?��\f
�^���8�w��U�U�07�:��=����h���K��Ǳ!�.�C���&����N!�`�(i3���$A�)�]eT��:
1���ƌ�j6"f���*��� S�n�(�a�&�0��eI!�`�(i3����,��=7�7K�P�l[�Ƶ�	���QC�Ҷ����S���Cu�;�R��3��m���d�0/0`9N1��-����!�`�(i3�,�B���{
Biۧ˺�s�˭;{o��n�(Z�ɽ��:^E��߆�p�hب�������kO�d��-��!g��J�s��F�e{iʖ.� �9�!�!*��*8����U[���*1tSjv���+�t2�;�������w�`L���JeJ��5�W��@�A٪�o�_&�
�:qEpj�E}4ظ����Ut�;!��Q�R��3���:
1����/�%�� ;̬gVdxQ,g�G��0��g�F��6M?��y�!�`�(i3��3�Z�#aȮ۔��5��Y��s����������,M끜�}Dq�f������!�`�(i3U�07�:�tMɶ���74/����G🕾{!�`�(i3�5ߧE4��ݓ�W����v��\1\����7��XW�G�<���>e)Յ�N��
�ge[I�/��kOT�H����g�G��0��'���C&8k��.ͥ�H�RtV�^�D�����0	�+G�c��=����h� 8�2�~S�e>%������w�w:�!�`�(i3��3�Z�#aȮ۔��5��Y��s��������2�(��W Ǳ0���%>�rGO�D mWNG�&ց�*�s����������,M�&U�)j�S��#�a�ĄS�n�(�a�:91�7��';��#j�ݚ�Н��o�t��8c���L���f�\%�F�w�[ޜ�}Dq�f��-�����j��&��!�`�(i3n��뾦�!�`�(i31���~��+�t2�;�������w�`L���JeJ��5�W��@�A٪�o�_&�!�`�(i3#l'U:�g[-�¾L���I����~u/��kOTfĉ>99��A0ok��(*�O�qe��0�U������KHN��R���
�Ŏ����ܐ�}��B7�Q�X��R�\��eN�q�Mf��=�@V{Z
�w�+��rdM�v���r��N�����?�d���&���n4s1մ�n:�z�'0l�L��������$*<!�F��66����~ω(�$V�y�2�x�h������M�!�y:i������M��j �M1����JV��GB%p�  �fAany�h�t��4����)\=��A���i9���Qp�	d��2������<�bሻ�״:��JV��GB%p�  �fAao�F)���;4����)\�uv�>u��d���!id=��¾ȼދ�Y"�I�,��u�C���L�s�ޘR�7h�,b0V�u�Q�ݚ�Н�b��
ߎ� n2ϒ�ȡ�&Y��V��G8T�w�nf�?ǉ�=�e�MW������L���	)��\R�][[�!�`�(i3�#�l+��B@
��B��+ H��*�{6��=��?��P�Y�6��!=.�
kZ)� [��v���Q:�7-mł(��gR� �ұf�?ǉ�=�;�.A�ى1�#��d_!�`�(i3�a\;V@|ऩ�jU/�\���WO+�jqh&Σ�h��I�
C���m�o��vPD��<!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3<�6�Q=�xsˁ�#2\z���L�f�\c`���6	D��&8�,�e'M�)�p��dHj�m�!�`�(i3m3�țZ��_�`I� B�!�`�(i3�<��N�Lf�?ǉ�=�$�V��bst�N���!�`�(i3�#ŪS�������k+#2\z��}�� �с�!�`�(i3�&8�,�e*���	�A�XF�����?UT>��˳����:=,3�/�r^�h!O���!�`�(i3frw��?�̞��>��vbëdP��_Ӯ\8�����$	�_:iO�A��*/�|��&8�,�H*W��u�a�ݚ�Н��>�@�C5]�꼧5#b|���Mk S���zǣ©���u��4��#�N�X�!�`�(i3�M����	�ĝ*"H�ݣ|Õd+�F�x�4zAo���E�{")8�*I]{�]!c�ߙҀL���Gk��,�:�N�*�x��0���>�	A�/ї:czZ�����
�%��!�`�(i3�����H1#�@;w�$C,0�?���v�h̤�Vl����S�Z;"�|q؉COt��t'�ݚ�Н�4?s����k�X;p`�(�����������	A�/ї:czZ������=��e��!�`�(i3���ٜ�]��/ӳxI�؉P9�?|�i�YɎ�#���?\a��4�$�~c/`L����D:f�?ǉ�=�Y=�Б�-��v�-���w:�4Rʹs=h���J	�J�y��*?(F`���G���}D���ݚ�Н���JתMܥ�X;p`��8
�[���oGt�Y?�Ɏ�#���?�5q{! lczZ����P(�s2�Q0�L@]HSϣN�}	E�!�`�(i3�$�~c/���Zs����Fz���oww��X;p`��5�j�))��<���wC������Ui�&xp�'��L���H��̣��h��N�M��� �{j��T7��v��w�K�B��f��0z�hq֤�eS�rK�
���ދy�'{w#/ B!�`�(i3!�`�(i3!�`�(i3z5:6�v�c�0T��~6j�"Hsg�2qqTS}ث�DȲ�w�ݚ�Н�!�`�(i3!�`�(i3!�`�(i3��n:�z�7�z����e�q�8��#+��
�Y8q�a~�'�� 7��
�+�0$��b��{��2������<�b��T5V+� e8�~��`��9C��Y�5��|��c���˫B�v%啖l�E��,��B�_��BL��N�]gR� �ұ+s�Di�R{{���5�&�q0\&���5��|��J�,B�v%啖l�S&�ɫr�?�d���&��ݚ�Н�!�`�(i3!�`�(i3m�ڨ�hծ���8-|�D��*CTR��ekl������a�h&t�iZ]XF�hx��G��!�`�(i3��D��������m#p�W��	]�	M$E�Z�ݚ�Н�*��^�"~H�𕎭own�~]�g����A��`-��'T���+��PJU��ĤI�v�����&8�,�e'M�)�p�`�Kg�'k�όz#�<Փu3v��U�DnK�]_!C6%K�pıy3�֩�U2P
�{���ݚ�Н��o�f�Ԝe���b�!�`�(i3�(�;\��B�}�� h9�}`A�)X�����(^ ��ߕ��`UNP�!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3�� л��B��dX:��+�k_����Zv���;-����`�����cm��x��{#2\z��o t�J�PM�Y��G%�&8�,�H*W��u�a�ݚ�Н��^yE⛀B��+ H!�`�(i3ˮF���t�F+������X:��+�i�	��_�V!�`�(i3-���
�I�>y��C��jћ@�/ʜn��C�(!�����Yk��s���eZ�c]��E���!�`�(i3Q)��Zl���w���4Wt#v���'w�?X}Ax���x��~iM5/�S3 <-���w�E�V{�!�`�(i36�R�W� W��|E�q��w\F��<��N�Lf�?ǉ�=%Y3(�6��B�r��!�`�(i3��l �� A����;���C#����d�E����'m�|g�~p!ۓ�ݚ�Н�&�2�������ȍry��	��b~y� ��&8�,��Om�"���^��r�VU���l����S4�0 L?�p���@Z����
� �!�`�(i3B��亁���&�%���B�'��a�[<�!��Tl�������l6��Q9���ۗ&8�,�cop ���6�G|��2��}����a#�fS��I���i9>���Ef�?ǉ�=�e�MW���^�yO�j���H�D���dݮ%*!�`�(i3���_͏���/ӳx��d��]�Q��f�_���u����g�&�0m����#oMS����6s
�:qEp0���Y$�8�$��`��7dh�?8X�˞�DG�e�MW��T��b9���ey�E�����$���f�?ǉ�=�#�m�-��Vi� �Znj��TAn�OZ@��5�h�ʪ%��18�$��`��UB�L5wG�!�`�(i3�:5A��p]M�|jHX{�t����՜�%P^���H> ��9�/�q#a�_�`�ю��x�T��ۇ�Qv�)�ˌ��Pg<\uu�����r����!�`�(i3!�`�(i3!�`�(i3�z_n�ԁi ���=��?�d���&���d.q��=�0��!�`�(i3!�`�(i3!�`�(i3m�ڨ�hծ����,�ǰ�6�Pr�|;G�R��Nr�",���ڜ��܍,6��zU�Ѝf�]P���Vr���J��:����p�m~|�֪GђP�#��r����2JHn��z�s�Đ��Xh�hk����`1 ���"_��̉�&�4C���=��?���D��ܒ",���6��*�x;��Ʒ&��;{ĥ�n4s1��>�w�Y�#�����B�@o��[�.r-����G��}n����ϸ��#|S������3[�u8�GLa���mdЧ^{�j-����h��t���oޯ!�`�(i3��I�Ūe�E7.�Z�"�4��%�;��7���ө�Rxem_�$n����������������i�^�=���p��R�f�?ǉ�=�w�Ylj;!k�2Nc��Nn%{�oꠓόz#�<���X�u��
)\Y��!�`�(i3
)c?�%Q/�}| �e����kn4@Q�/��ݚ�Н����S�|J�X;p`�B��C8�4`�Z�l{?V��j�c�[N�&ѐczZ�����ݫ&�b%%f�?ǉ�=��=m緒6����}F��(ja]p�X�o|30��^?8�$��`���	(��7��P�v	��Y�Q9���ۗ&8�,�cop ���6�G|�</Sn��-�¾L��S��I����yP2Ni�~�ݚ�Н�*��^�"~H��
�[�<�`A��_i¼\K��
�:qEp0���Y$�8�$��`��7dh�?f�?ǉ�=�*46;�[-��$ϙRl�bu�	?�cx�3Lv	̅��!�`�(i3>N0Θ��ݚ�Н�Gظ0�����X;p`�l.�	�C�
�:qEp�����%������r��	��
�Q�}��"���l<o�;)�y�y������x���m[3�� ��
m}:[�O9UNTnF�\F�l9Z��b�Bϱ�\��FHѽ����8H���&�bP����|�J�=��?R�����!hh����P.���ݚ�Н�!�`�(i3!�`�(i3!�`�(i3��kw�G��.�g3Zꢯ�wv��ޟ��}tt��wN�p%
-bK��:z6�U���e����T�bC�9/���U��)���Y;e�iK-pm!9�>��n4s1�U��B��-_S���\���&�vf��G���"sS<GYqcHTX�';��#jx��7��� �ؼ��"ª���!��"� +}0�ʂ�j�Ï��	�l�lM�3 H�RtV�^g�G��0��}�m�'�M �cJ$���hpI�_�c�r%�[�ap�Vȓ�"����Y�5ߧE4��Fr��j�p���"k��yV�:���(�'���:?���