{# include('templates/info.v') #}
// NABPMapper
//     3 Jan 2012
// Provides addresses of the mapped projection line for line buffer
// Outputs available in 2 cycles
// TODO reduce look-up table size by using symmetry

{# 
    from pynabp.conf import conf
    from pynabp.enums import mapper_states
    from pynabp.utils import xfrange, dec_repr
    from pynabp.fixed_point_arith import FixedPoint

    a_len = conf()['kAngleLength']
    accu_part_fixed = conf()['tLUTMapAccuPart']
    accu_base_fixed = conf()['tMapAccuBase']
    mp_accu_part_fixed = conf()['tMapAccuPart']
    mp_accu_part_shift = mp_accu_part_fixed.fractional_width - \
            accu_part_fixed.fractional_width
#}
`define kAngleLength {# a_len #}

module NABPMapperLUT
(
    // global signals
    input wire clk,
    // inputs from mapper
    input wire [`kAngleLength-1:0] mp_angle,
    // outputs to mapper
    // mp_accu_part {# str(mp_accu_part_fixed) #}
    output wire {# mp_accu_part_fixed.verilog_decl() #} mp_accu_part,
    // mp_accu_base {# str(accu_base_fixed) #}
    output reg {# accu_base_fixed.verilog_decl() #} mp_accu_base
);

reg {# accu_part_fixed.verilog_decl() #} accu_part;
assign mp_accu_part = {accu_part, {# dec_repr(0, mp_accu_part_shift) #}};

always @(posedge clk)
begin
    {# set_eat_blanklines(True) #}
    case (mp_angle)
        {% for idx, angle in enumerate(
                xfrange(0, 180, conf()['projection_angle_step'])) %}
        {# dec_repr(angle, a_len) #}:
        begin
            {#
                accu_part_val = conf()['lutMapAccuPart'][idx]
                accu_base_val = conf()['lutMapAccuBase'][idx]
            #}
            // {# accu_part_val #}
            accu_part <= {# accu_part_fixed.verilog_repr(accu_part_val) #};
            // {# accu_base_val #}
            mp_accu_base <= {# accu_base_fixed.verilog_repr(accu_base_val) #};
        end
        {% end %}
    endcase
    {# set_eat_blanklines(False) #}
end

endmodule
