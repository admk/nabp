��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-K�趹���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�s8�R�	��q5.A��|�H����VM.H�{�|�w8�M�Q�"�,�#ѷ���� �\_I+ĂiW,���D�+y_�L_H��-..i=?�m��+�<4��ˌ��|��v��ӳ��$Fe@���N�w	*D���y&�f��+K��[y��ڂ�1aY���~a1k��1�/lt�3� P�;��1�-���f񻲗��~o��:���F�q�\�7Y[���G���d�֗r�5�c$e
�9��Ax!P�������H3����^�CG�1 T�V	�tL��	�<�A�}Q��	����<5�T7y;��S���4B�@T�,�찱�y�Zk���fi���60��g��b#Ӡe��?�F��&k�ZV"��s��;#�A�v�N<��;���u��w)�S�5� ��~篟|�<8�F�-:��ԧN��78�:r&@��$�9��_,n׎ ��73��>g�����Mp᫼���hvK+�va��2鍔�	g\A���V�2���y�͌�4r�O��C��0���df�����_0�M(5>��u���;�Թ!o�o,%H�%�ì���Tl�
� �AH�}��� ��fD���N�J��R���S�!�� l��F@�4%��%dZ&��Ǯ"�lf�~��m���w>�K�6���	x]́��D�Q���X��� L��57�8O �L#���O[���StI��B6:�4V�f��n�GE�y8|�g��P.!܃��L~΄gO�3�q$��nK� w�;�d���N�tכ݁=9�|Z���ߐ'�[�Z���1VU���+L��h��X�vB#|y{����P7�.yt�gU*Z9B[�^������+�ͫUz����~2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcMD��y�sY2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc.�
͹U��|�#A�)�(F�ow^�\JO�F'���Xw��4�L�3�[���A6����ʌ�<���o�3t���!ʞ�b�F��?�Q�E��GW��e/?�s�m/C�N{a�9O!JoE'U�Y�y��
r�)�Y¹w����i��T!ix�AH�k[�^��_�)��6�$`W�����%3?���kW���;��sD���L�S5H�j.F�H�J���E�L�Xڈ*-}|��ι%9��oGo�Z�J��ݪ�ufҷGپ_����b�[���F۰2�(����5��x���|�:S�Q�[����g��㙖s변�u��i����*�{¥������z�)
ԏ�.T٢ߡ[p40�zɈ:��B��J��H9'E�HG.���hm�F!�`�(i3���P!�&K�A�H����8DE��	�J�ILo�����,[$�	J���GKer�I�F�ݦh�z�(������l#��䩛���y��lD&خ.�o�O
��^O��w��ԩ9����'*D�]:�W�G����?+D���0�7a
��r�yد�9�����~���-�f�t�������~��(,R[#�(y�T%ME)��!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3o�kr�.z�o��x�v!�`�(i3!�`�(i3!�`�(i3!�`�(i3<�6�Q=ؿ�?��5Q�Ub���Ɩ���2�Q��0m �]vo/~�e6j���-M+�Ԝ�}Dq�f�!�`�(i3!�`�(i3!�`�(i3!�`�(i3zZk���?,�=k���52p�8s�?�������`F�k�d�l�!�`�(i3!�`�(i3!�`�(i3!�`�(i3(2��\YV6{,q3�+���C��n*�k`��ͯ�K����6��~�?Q!�`�(i3!�`�(i3!�`�(i3!�`�(i3_Q1������t?uw|`�ڛ�m��e����2��=!�������Mڂ+!�`�(i3!�`�(i3!�`�(i3!�`�(i3�1�?	/�V�8��/��6�?��h�0�����9��S]��ݚ�Н�:��9KmR�^Ƒ�Ӈ��t�9>yh��DvO���v"�N-�T�\3%/��.�@��RN�]�5'c`�/��ȍry��	�s�٩�삠k�bWbG@���p���ݚ�Н���?��[� �V8��v ʞ���
�:qEp� LTx%�0�أ�Mft�s� u�?D�8�镁�aR�!�`�(i3�i����u��N�v{���df"�	-7���C��L�c27���&�_��lC��U7�C��zC@��f��p�(p���	��
�Q�}"�4��m�S⏸[��]2�y��]�!��	Ǹ�y85��9�L�fG"j���b7Z�n��[��{_8�Y��=�}�Vݨ��}Dq�f�i�]ʺ�
ǳ��ٜ�]Ǧ�JS�cbp��'@
9��y��5�%]�����3�(���tP"7��%e��0�UX�Pp42JF��c;x�@Ã�D譸3L�*}F�x�����Z鎬����Ĺ#{����}Dq�f�)�{6�U���ea��L��K�*� ���G1��[��K�+EC�����6��lC��U7�C��zC@��f��p�(p���	��
�Q�}�d4�n�Yct_��צ��
t��{<���낌)P<�ܓ�Y���aR�!�`�(i3m����'K���Æ6�HaDl��+BY��9��8������{r��;�¬pX����B����qe�@Rv���|z�ä�@��m�r�����I���`��`�v����2y��l����4�n���xǊ�Jם��t&:���a��2��1�V����(��8fDs;ly��\%��'T���+��^�Y_Ez��!%���Kv���ft�s� uƍ2���lğMg$9�rJ
_�y�V( �w�;>cbp��'�����C��ݚ�Н��l��#�}��
�'����j��<ͧ�:|��b+}y[���S�fDV��,�����
�9�j���B]��>��y���|e"�7؛ڇ��lԇ�-{�(��̓i��:|[%.�|Tck�=�mJ�0�6��q�1Ig�I�?g�f�(�r���`�s��;#�A�vȹDc�c~Op�����M�v�j. �	(?��I�?g�f�(�r���`�s��;#�A�vȹDc�c~O����� (1Lô ��q��Xx+�~F�5�q��[4J&)�훪�K\����H� }��6Z.�m�$*���Q�q�v��+BY��9�?�>L���9�����x�����s����
mO�h��M�ns����V�Q�q�v��:�����`�@��i�&aD�4�Iv(1B�@���p���E�qA�y�=0��#���t{��*��f`��$^�����}�
�?��9/u�6��?��{�:2QYeƈ)P<�ܓ�Yb!��u�m����'KȞm�2GS��]�!��	Ǹ�y85�5�_k�XЩ�c��><�$��W��_�ړ8���/�l|�*"k���(ӈ��Bm���8�� �?,MU��%�kˣ����aU)`k�]�!��	Ǹ�y85��3}�@�7"j���b7Z�n��[��{_8�Y��=�}�VݨC=2崝�g��gQ��(鍏��pb>$y6s��&��J�C.W26K�~��@���Jٯ�n
�5����`K�ӄ�B�Z��a\Y����+���LQ��a�\����BP�-u�"�̞��>����-M+��*������:������m�5��C�F��$�ilG 9a�{���B�D�F �h�`�>��򴏓�	�^4�:U�>��Oއ�?t},�׉é]���k��S܇���+�]l�B�:	�.E`B��e��Oއ�?t�<�VV�$��
��:d�z��ſ��D�d
 � v�)��& �8�C]H���L@�B�_	�Ƽ�E�����H���L@�B�&�(���D��)����>�qpNɡ���t⣟ڇ��>j��K�ݚ�Н�B7lĺA����B^-#���#5)�!�'dT8�,6�x1�~g_�	y�b�� �S3�
��G�&���\�<D�!�`�(i3��<㡧����5n'�	�4�_��2������|�Y,a�/̆��B0F�z"f�ú��g�=�?�S��O����R=l�ֿ7�8���ݚ�Н�!�`�(i3!�`�(i3!�`�(i3!�`�(i3"�9ŭ,�]g�tҬA�E'�ТoT��!�`�(i3!�`�(i3!�`�(i3!�`�(i3���y��lD�X6�4��Ʀ+���(9��&s��<�9��W0��!�`�(i3!�`�(i3!�`�(i3!�`�(i3<�6�Q==d�Ɇ�;c8DL���7��){�%��!�7qp��k)!������f���	��+*9x���С$�)�vx��?w=�B�ht�&H��߷~��nJ!-ȹ���1L��	�Z�kfc�_	�Ƽ�E��������`+iYbx{^4��*m!�`�(i3'E>�����Y��a��u�k�?.;u.'��3&5L��$
c˃��o���G�ب:�T�t�74/����L	k���R��UB�n�5ߧE4��\E�W��4b!2�͞nOYw�,>�e����%�����C�^�n��3�t�z��z��_n���-�+YF�����n4s1���=����t�n�𤠊ջ^B�}u��ݓ�W������WS�;�r��q+s��J���ƍ2���lğMg$9�r;��`�x��Υ�h�B���|e"t�td���5��Aڬ&W�\��.��4�zm�$�ܻ�u��r�����S�f������f���ݤu��!�`�(i31���~��'T���+�N_��ʥ�L�H�l��ݚ�Н����F��O�/�"����03�gea\�3��Y$��s-e�Z&��"��ӌ�r���S�fDV��,���S�i<���%��Y�;�jmT�#�#M�#/g�zm�$�ܻ�u��r�����S�f������f�=&`�G��}Dq�f������!�`�(i36Gި���74/���
8�	3�fĉ>99��j���GpG�&ց�*�&��j���3��Y$�1���/������E�EqLt��.fĉ>99��|��3��׹�>d���9�eW5�2]k�WM��q�U��)��G0cE��e`�:�N���O��h�U��B��-�Q���Q�@}Z��u/�M��Ε�`UNP��D#�]�q2&U�)j�S��UՄ��g&xdp�؜�}Dq�f�,��e�R��	����;�jmT�#�Ȑ�TA��M?��y�!�`�(i3�L	k���Y��[�P@�m�T�	��x��ݚ�Н�z��SͲ����E�EczUEg�>fĉ>99��A0ok�ݗƩ�2Z�i��/7@Ã�D譸o�;�6���|e"�#M�#/g�n��뾦��mJ�0�6��H����Yq���3������&G�B�'��a�]l�B�:	74/���
8�	3���w�w:�!�`�(i3�L	k���Y�٧�i_���HN��R���O>�R�`m�ڨ�hծ���'��@�my$�N�z��SͲ����E�EqLt��.����1��b�i"���φ��<�6�����VR�����_h���3�"�l���k�b^ � v�)��& �8�C]H���L@�B���5Z2URK�a��R#���`+iYb�����&G����ł��cЉ�M��˿�񴞻�(ӈ���m�r����:#�R_��L���;^�'DV���b�z'hۉ)��d�7�q�o��w��6_�۰��ݟ����)�Y���4#��Z ���>6;��'j v���)��_�mS8<�n������_���s	 j��̇��'_���s	 jQ�F �:#�R_��L���;^d������`�v��,ƴ��o�;�P�t�5���F��O��z~S�����U�_��ȧ[�դ�K��R&��	�|r>�ei��F���4 >y�;o�� ��'*�ha�u?��F�zw�^��S�&�2�"G����4 >y���H�`m�6i��̨D�'bʟ0�}��'[�M��)��c�X`��_/�.����d7����wo�͑A=r��ր��z�)�._�g����+�ϊS �i��{�I���;E�@Nz�?*��K��Y�R,���]x��� ��W�҇��TM��o�u�/<�KǣDy)ʩ�3瀽ݻe쒮�Wf��K�4~FD�fT�wRyAx��PS�_ ����/�XD���^T,[O�5�:1�x�<b�y��tqӑ�l�n�ZlӜ�g�PUrӡbZ����YaD_A���f�Ԟ-zq4�0��<�\Ys|��t�Q湟F�-��1�,�� ���BG�
�\ɦ;��|B <�Az��S⏸[�nF�����2�[Q "M&��?�d���&�R����LgHE�$�N�P��(�3�.����]9�(b���*5�����e{"�Lެ�k�� �����=y����Y��E�
_���s	 j'��|@8q�a\Y���R�^Ƒ����"X��[B��r^�Z���v.7a
��r�H��=q�� �r���җ6j�"Hs�u����$�|����ٞ}aBVG����8�3�M)p�ۉ��?�d���&��6)��Tj�`����nK7͍��ճ��)��{��&^�E�6��������`:tUx��C}�>��$�t?�@@���ތ��t�h�y �R�r��̗{�4���+�".��cЉ�MRbv��[{u7a
��r�"j���b7R��~�<��V��	��y℺�>��3��0���藘�������7���