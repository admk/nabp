��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-K�趹���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�*���g S��/P�p��]P*m�x�t���E�L#uc��WŬ�+�-ޗ(huUPy�����h���!�}�1�:�Ω�*���g S��/P�p��]P*m����)O��Ξ4�"�\�� ���K�O�{��
2�D��Sm�f���=c\֣�I��B���t��|U|�/֚m� �+d��.8%D.��n�P��<�!Q������Ś��
��H,7���ZXWL�sZ�	!w���� �bRw�����IL�+�{Dr[��:�\��~���"��y0��9�QH��������\҂�% B]�pE(���B��|�o�r� ��J��ݪ�ufҷGپ_7\F���r��RL�a)ѻtUWR��]��5t��^���Y���t�&�7C��Hl�>7��yx_/�Z�s�	�=5�NUD60L�U<���;�e��e����[�/��2r�O��C��0���df���z�!%���`�򾄖�u���;�����6�b'1�}��)��gi�HF��eUٻo���mi��*	�ť�.^�i��' 1wH�x�xs��3�<A��z����
a�������~�+��,/,����W >g1�]l�&Y��F}갨y�����# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��`y��f2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�����g��~�X�x��S|�m����Y�{'%s#K�v]|nf<�,=K�F��N��j��D���s�촜g1��rN�.[4<�6�ۉ���2=�l���������Q���p��^2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc:#�c>�ϜT��:�E�>�5�4W�g`%J��N�9��N�^#?���E:�J�k �?!R��	k�9ːh���%��A�뱛+ƯE1j$,�����������ӯ������@	�J��l-[�v:v��M�H
�}ʊI�٦�D�`F��al����Fv��ߑ9��E|+�5�(�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��T|ރ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc{�-���(��#��w��Q<���2� m��J@BY�?EW�j����qS���+�>����KiҽԺh:�jޒ0� 	��F��=?��m��&+�!nZ�!
���>X�J H��K�zk�����x<E����^��%S��I�JT����Fz��l9�ղa_��=J�^���,��͹o��Ca2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}�߼
�dX^�	9�e�Ч4m�C�tT��A��蠿����d�Uf�.`�Z������"��y�R���1x�]�^�[��n��iܕ����������a�"�5F:	��,&�<3Ϲ%�o�ċ����q�ʈ2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc؆-�qh��7&n-Ȅ�W��i�4�Q<���2� m��J@BY�?EW�j����qS���+�>����Kiҽ�������.�񈉝��s5l��o�A
��_�b��Xw�?�b�>��O}��H�'1�w�z���vL�vO�
�rU�?���?i����k��u�� ���$����t֬s�'2�o����"�RS.�E!2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>hN>�4�
��C�<w��>�8���Ę-ai.���@��8���i�E̳&k	�I]����o��Ca2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�U���2��-���MV����U��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��T|ރ��Sc�j H�g2��\�b�#��lWY��lz�M{�C��aO/����N4Ҩ,Ű����!d�h��<�q��7܌:���ġC����F*D@��j�5�a��3Ն��ج5S�ޗ)�t�!�Zu�����@
H$��jg��+˘\5;ԉR���F����!d�L�~��&����/�5�f'?	G݈�����a�"�є��E�t3�Y	���R���:K�-�D#q��4%G_��-���`�r�e��\
�z�.��a�S.l"�%iq	�g���H�^A02�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�JW�_N���4ҢB�'�;5�3�����љ2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc���.��(�Ze�eu+�1Ƙ���<�<Չ��
u_�^�6Lz�#j���ؾz<�hjݭ�F���E���%�a���b<�d�w;��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc:#�c>��`ݙ:���߼
�d���D���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc{�-�������:�3y�Ƕ�F������G��-͕��O�"�FWy���l��s1p��"nq���z_�3���4�듴,`Y�{'%sa�6���� <&�M#'���Xw����s�c�"nq���z_�3����DƯu&7���F�!�� <&�M#'���Xw�h\K�5~���:�3y%r��QuP�T�UX��v�^ܯ�~����pؖ-�/�+T���u�I��U��؀N�&jl��� Ϳ�$��0z�cUL�|��q�A��R� V�pό���.�N>�4�
��+EmI��1� ��5}�Yq��T��h��<�q��7܌:���ġC��חsܢ�2�����"��p�~ �����D��v�j�_���\'?2n2��;���!ocN�RZ�N�X�;LdG%윈[R*$�s�,�TMo������a�"�_����h�&6B���U���e[�.��<PM�Q�����-�s�<���dL�t+�R�+���O�AJ�㗲F�hݿ��KD�[R*$�s�,�TMo������a�"�_����h�&6B���RdM�5����$�(�+�j"i"��L�a�1!�ӯ.�����iM0�3g����ޔӺ�(,��AԢ�a\�w�?�b�>޼�\�vũh\K�5~�#*�F�E�����]6�l�(�3�i��%єX�S�EP"G�wk��a�S.l"�����x�W<1i��|���F �������X�c��z��^���m������"��yu��������DƯu&7���F�!��t��\����b~�ff1�^����!�']5����P�;߼
�d4I�<w��Z�^T-a�ؕJ�w�?�b�>޼�\�v����T�Ŭ��j�P�tCu^(򎍖=bT-a�ؕJ��d�nX�RM��A���va�{���ȳ�I!��;�Ɛ����8��x`��������D���J7"��10�����S�����H�
B#�ۉ���2=�l����FqqDt����D���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h9��)�N6mj�N?����;t>
�o��Ca2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}�߼
�dX^�	9�e�Ч4m�C�tT��A��蠿����d�Uf�揆0�бԧ2N��n���?���^��a�\����Nf[8��(&�L���p�`�6��Qu���% gWVbT+xΣ�}��Q?M8�f2���u�䯄���\�˺�KA2���ݚ�Н�
ҭ�3���]_�t?	�$f��_Ub��7��G_��Ct�w#��@������37y�����:���b��qeҽ.��>���Kp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 �_d�Jq/W��������f�o'
���#�l�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcT���u�I]�I�rT�8���|�F��\��:���Ԑ���e����޳[��g6�w�9\S�HE�N}�m��{B���T�Dʆ�In��t�8&���I���|I���a۲5�����}Y��	}�@��O�׽����Yk���~�	�0݂S����B� �b�З/��@��2C��'� W>���������F��O�}�	76�&�R�Q���~��p����B�b�>JrP����p�(�6k�4d!��-}�	76�&��A0ok�����a�"�_���3� �d��f~vW4��`��H�^A02�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��������Q�MHf�o'
���#�l�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcI>����a�AJ�㗲F"Wm��|������
��s�����E���%�a��s������XP��~�26��\�o�mW���5F:	����n4s1�ЂDa��(�_�R�G��=�gw�⽒��Շ9�/�|#HK��ehj�t��{r���B� �b�З/��@��Q�����;b�-�2��;�P�t�5���W0�]��e|)0����)�x���3�}@��9�ڮWqUv �6U���Lt�{��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 ��M(?^v�,�mI�p��o��Ca2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcT���u�I7.���K��r�e��\
�z�.��a�S.l"�S�)37J*u�1��r�p?��$�Qu�&�<��G��d�٣�����c����յ[+8�
ҭ�3����h��]�z�[�+�߶37y������(�;-�(�ь�$�5ǁ�O2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��T|ރ�V��݀�p�5UˉB۬�o�W`���s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}�߼
�d��f�u�q^����:�t1�$8L�~��&�a�'�%~I��U�;��r O��M�Zb.�Z����$�Qu�&�<��G�ȵ�ixUS�!ih���S��T�\ �͜����Ƀ(����<mlXw�X�*xlL��I+=5�zߴ�� h�ҩ�N�D��泵~��zq����1����z�F��+���n�)7�h��T؁��D393�5�a��3�tץ���:Z{G�i�e�n�^���Ě�����Qu���%��,�,
((���G��)��4���S�8B`��@(�6k�4d�#��M&sǚv�j�����{]F"HN��R���מu��� �H�0��
�U���G��&��/Q�g��U-�ex�����">_X�;P��ĆjS�O��b��֔l3��$!��qR7׷�:�Kp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h���\���f�o'
�Us�6�И2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��AX��-���`�r�e��\
���F�!�� <&�M#<.�_&|"�ֱ�q������m�q�C��l"�u�ȅ�Yt��1��IM����`y�����n4s1�ЂDa��(
��B��]��Qe_%r~J�3
�$k��S��c�ط�¶�`�aT��3Gs   ��?2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 ���Y�Q��bz	>Xd�|!�x��02�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcI>����a}�QU���B+�0���a�\�������޳t���92 |ȟ���èVR�@�6�֐k ��J��?����2��<a|��tʪ�q�G��Q>�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc:#�c>��J����C�qҢ�����N[ m�N2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�o0��U����開���-P�ȳh�L>s�]�!��	Ǹ�y85�E���%�aS�)37J*u�1��r�p?��$�Qu�&�<��G��d�٣�����c����յ[+8�
ҭ�3������NM����i7N�_	�z�w.{��w�_��(�6k�4d�{j����}=!�ҳ�ϾQY�u��A�0���򴶽!�y�"�V��5M��z�o�>��U^�����v�/��xv�3���\��:��AԢ�a\�w�?�b�>��]�!��=���W�N}�m��{B���T�D�]�!��`��j(&�L�i��ko�$�?D�8��R'cf����T�x��QU���^4��y��j��kL1���oBΒ���PW!�w(�y?�?�JY�)�֬w�J%�H���3�}@��9�ڮW��Q>�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc:#�c>��l�W�z��Қ���lW"`oG&2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc\�BDL�c���w?�����XR�[R*$�s�,�TMo������a�"Z鎬����Y8�Sv�~�26��\�o�mW��Z鎬����+�E/(��^��f��-)a��m5i��"`,9�H�Wq�71�ҁ�\�$k�Xit֭�h��O��W�	Ⓤ��5$r�t�}iCt�w#��@��S��c��څH�8��)B�>T���u�I��U��؀N�&jl��� Ϳ�$��0z�cUL�|��q�A��R� V�pFr����A"�U���w�c*����W"��ό���.�d=��¾ȼƸv��*Qxm�QA�Q* 5�����}Y�]��h@�YyZ��}�Q?M8�f2$ Hl�]���P��))O���w�_fHN��R��Gu�"�0�R�@�6�֐����o��4q�I�w�o2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc:#�c>��kB�1L�|� ѹ�8w��4.\�����s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��T|ރ���-��ԣ����/�ʹ�z�$�W�@��!���~Pw-�h��R6ti�7���x-�t(�Cy�H�Ek 3��㶺���cJ��e�e�s.��"���N3����k��!gp'&��ͦ	2x����$˾�T���u�I��:��l&�!�Ť̚��DƯu&7���F�!�_(����@҄���G��b�i0[�S�T"�IÉ��,�,
((�H*�iH��[��(����Aڬ&W���O��G	_�mS8<�n�ݚ�Н������a�"]_�t?	�$f��_Ub��7��G_��Ct�w#��@��S��c��Ny�^YC&��Y�g�f�����s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}��_�����l�!�%rf�c�R��kBޫKp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h��g�jZ����"��p�~ ����#V�&�t��c''����:�ui���?8���yB-��fx���{�h�)ȗ�bB˶s.RO�#C�R_Ax�.��Cɹ��e�P�~V�t ��7[�ck�?4�V�ʄ�Z��AJ�㗲F�hݿ��KD�[R*$�s�,�TMo������a�"�'n�^0o]�B���[d�#��Ӏ�`,9�H�Wq جI��A����� ���	�|���H����y(U���������u��r��ʥ�nr]uxp=�*.o�;b�-�2��;�P�t�5���W0�]��x@��6�����-�������V1�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc:#�c>���Yq�s��Dn�k~3
�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vch��\��f��RdM�5����$�(�+�~����p�5�Y�w����9�<���N>�4�
����(�.P�3XRt%3�o2C�g�kgw�"��I66�v��G���V>�R<�2N��n�O#H��Ek�x�ZWEב.`�Z�����èV��NƥN���˟y7�%M��أͽgF"?�nק���۠$/I��A���Yk�����)g��I�߷�c/�B� �b�ПB�'��a����omi7xob.�Y�2W>���������F��O�}�	76�&�R�V�"�0ɶ37y�����=$�B�>�o��Ca2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc%�d��x�d�j]�\�2���`���|!�x��02�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcI>����a\�����8P��=.���\��:��AԢ�a\�w�?�b�>�P"G�wk�8%PT��&��~�26��\�o�mW��AԢ�a\�O7z��4�dQ-gtյ[+8��i7N�_	�z�w.{��w�_��(�6k�4d�#��M&sǚv�j�WS˓C�^��@�VҒm�fF�5.]������������^��x��/z*x�n�H�^A02�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc{�-�����J��zI�R��kBޫKp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>hN>�4�
��3���<pb�*(%���AԢ�a\�3�g
�!���U{�:�E2�,���I!�`�(i3!�`�(i3wi����C>�F��}��T�\ ��L9�{m��$��$�Qu�&�<��G�xZ��j�
��઴y��R�e�0��|#9���W>	����h5�����}Y�]��h@�YyZ��}�Q?M8�f2౉+�+�����>M6H�O���w�_fHN��R��Gu�"�0�R�@�6�֐[�%�g��pl�4ʀ�$��B?V����s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}�ڎ̞i�6����������R��kBޫKp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>hN>�4�
����7��M�&\})������u*K6H8!��vp�P}��O��ꅽ52����$�Qu�&�<��G�JHn��z��
�kˤ��.��|ȃ��X%)�j�=�|�86� h�ҩ�
ҭ�3���qՎ0�W䪸�M����'{w#/ B$ Hl�]��J� s�HN��R��bP�63Z�t"�Ԉ�F�Ǎ��ݸ���g�b�?�D"���Vbe��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc
MH���ﱾ#c�~�����@�_32�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 ����"��y�S��?��L�����@B])�+T�b9���M��A���va�{����PD}#��ůN}�m��{B���T�D��\�v����S��5���n4s1��7�癆cg�>@����7Bˡ����Y�y��j��kL1���oB�ԝy'����F��O���S��c��څH�8��)�rs�U��!_S�~��p������8<�V�Zs˿�}w��ix�AH�k[�^��_
�o����L