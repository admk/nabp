��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-K�趹���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω��:%��Z���xN��g�.H�{�|�w8�M�Q�"�,�#ѷ���� �\_I+ĂiW,���D�+y[ف���rn��mo����/~.)��3�(����C�X��2�k(����)O��Ξ4�"�\�� ���K�O�{��
2�D��Sm�f���=c\֣�I��B���t��|U|�/֚m� �+d��.8%D.��n�P��<2�q�U��k�8u[\E���@N1�w�0XL����[fe�Hs��9lSUQ�S��)���2Ee�Y�R2
�I.��	���
����k�������0�?�}4��ѕ�������U��=>bMab�	;4��G����a�����(�I�?g�f�k%URPx�ζmR{z�W ���������	x]�fX�eϝ(�Я�mڍ'T����X�w{������:�%�+T%2q򋙔�M-US-�8<�n�У�Ǝ!�ѠV�>!�/�7��u���nEA?��m��3t��⫓���RL�a)�ƞ��U<Bg�3���M Ce=6�([a�EF��7C��Hwɶ R�p��4�s4�o�qR��p������M<D�7�s)	w�N\`�a���!4d���-sk �0%̄sb�� bL�k>F�泂�0�V�@���RL�a)ѻtUWR����H7��7�ޑ����<��&g�7C��H��C=�)3�C����")�E�'3H��[e)�p�R\��ꫜp&C����/B!,�G�;(�B�T0�z$�}���E6sC&�gG��Hc�e$���=M��8�w'��(�D�&�〨����cZ	�M2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��~ǳ�!2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�tw:g�V|�hi��p�7��Z鎬�����R�LM��ħƿ�9c�5(��}���SaB:r���q P�^�&d�A|�1�:�Ω��]��
��rE���ƪ�(����D�I�?g�f{ì(Q[nS5H�j.F�H�J���EJ����%@����BF+�va��2鍔�	g\AufҷGپ_�	g�yߓ����<�m��+��$|��;D���J7"�x$�^w��aC�h�>�N{a�9O��Yk"1/]���!E���VG%��m�q�,�,\ަ�It�k\,آ()���;��G���9��'n�^0o_
-��[�����Kp&�@���k��l0��F��jT�����Nb�?49�����_�\G��4�	B45k�c��`��'n�^0o�!���!��x�	�2��g�P�e�9�:�]�^��'n�^0oM�D�;��-+0�l�R<�q��f�}��Gظ0���������5	���]���>����C�h�'f R�����5	���]���>����Cοƿ�d��������5	���]���>����C�?KYC'v�������|g�Y�'���Xw s4S�'�i��`�z&"hkIH*���>RTت�I7��-5��6��	���`y����ꢤ�Og�[N�&ѐ��(�
t��Y�{'%s���'���ը��_�\G��4�	B45��lC��U�T�\ ��Tǯ�!�tӱ1R�m��+ r���7���?�_���>3��w-iu�`���`�+N��?���&���#�{�0;�}����\Ҥ�Yk"1/]���!E���VG%��m�q�,@���j|Z�a�P�Fpwe�2l��4�y��ɦ�@^7&ģM�'n�^0o�<:�W�_ĵn(���˧�0z�cULjaGkƊ~F˯�+)�"j���b7|#9���b!��u��<��>�ڍP:�_?�ia�P�Fpwe�2l��4��a��se�ξ���X��9cѶ��i�ܰA����sC���"��|����{��$gOv��Ψ��F$��O�&��������v$��fP�'ׯ�߇&"hkIH*�=��#�-���w��l��ML�f���|����OxtX+�Y�8�>r&��0�~?5+�oz�oVa�x����0/�e��9�S;�¬pX��g��U-�e���b P5b11��m$��O�&��;�L���9��Xv7�j���0/ܤ�(g��VO�f�6u �q�t��},�׉é� Ei�lmZ/���@�ܡ"�,�>E����+����eǎd .8����*:W�q�ۻ�o
]�R'cf���³5��)���;��cj�-��?�d���&���5�G
m�tooS�c�{I���,'�*;kO��u��<��>�ڱ���
# ���0/�e��9�S*V�M��nD��;_��8W�w��fD�;�����Ǣ���ϜB?�<&���}�����z��i��xl+r���y�����aHu�4?�d���&�V��o5]���aU/�`,9�H�Wu�Σ�����]�8��r�`�c����{�v�$?�d���&�������y�F_���ٱ'W�w��fDfTYQ0b| ��%UG���.J7h�_ݑ���J�󈷛�'�2�w�0�9�]�8��r�`�c���ՍPhT����Z��!�`�(i37�! ���]�IX0F�MV�ҁGG�.Mm-;�!�`�(i3{y����:�*" �`�H����Qw�c4~Nr_�mS8<�n�ݚ�Н�SƏw0��A��6��
��=<�6>e��0�U+�qbp@�!�`�(i3�k��^�1Aj��t�35L��$
8��2�ֈe�cN�0��ž�Ć�T���7X���c�}�����l��=�O�-v�*_�mS8<�n�ݚ�Н���'T���+�;�7��w�����$����hY-N�g� ���p[~3Ħ�0r�/)+?����7Ա�D��,H/��!�`�(i3�5ߧE4��!�`�(i3��Ě�����}Dq�f��Fr��j&���"�g7�}޴�z�I��)���W�w��fDA���ő��}Dq�f�Ip��u���v���$hk���@8��m�F�!�_H^R |~�($U*���yf��>5�O�%E#PZt%��m&<�!�a��T�o��_�Rv�䩲$���dS@Ɵ�o��6}���iI9�o��ݚ�Н����"sS<�0�zG�������&G!�`�(i3!q��V�ys��e�sb_X�XV�b�z'hۉ)��d�7�q�!�`�(i3�Ro�G/]%�z�-uͺ�s�η3G��Hb+�����;y��v��\���
^�ݚ�Н��H�����Yu�������&G!�`�(i3SƏw0��A��6��
�g�����;�7��w�@z�צ�:5A��p
�:qEp�;�P�t�5!�`�(i3���F��O��ݚ�Н��׹�V���$��b@��ʚ����.�g3Z�)V��B�1�F(� 2�}}�	76�&�;��|B�:[c�ϲ�[F+�t;��|Bm/�Bơu$m��{Ձ��cI�*(�'���Xw�j�7��\F��wG,���_�\G�k�y'��a`��Dq-/%�FX���v�\�b�U4��\w��˪?�-X��9cѶ�����ڀS��d���!i秭�B��@8GS��`�ƫ�P�A�I7��-55x|���MM
��,=?�d���&�t�{#	�x��_--���g{�C����c ,��rQ3���w�@V��t`x;��E�i�m}66j�"HsX�q&����*�HZ6j�"HsӋX�k0��7��D�)k��m6[��-�b�+�