��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-K�趹���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�=A���>�LZ*IV���^���������g�3�7x��������&�ǝ�+zA��]��~ا@H;�W ��W�5�k��O��ڴ���WЋ��I�?g�f�ja1�n�[�c�/�O��?�;��XC��o��y��b1Ø^���#K���lӧIA�a�V��R�5K�yQb�I��68�/�YJ�'�دv)h�V~�$v�p��"}�vo7k2a��pP.S��*����طǪ�`DY��YH\��!���1R�_ߥ�]��4�:j�l�,9��)'��e�Ni�H�f���Zߧl4���0�?�1~�x�c�	�L}���i�m���w�*��O0�To��6�*�2���K{l�+ ���M�� ���M��z�Ft�f ���M��z�Ft�fz�Ft�f ����γO���Fz��z���y!�`�(i3�z���y!�`�(i3�z���y!�`�(i3��Ͱ�N�ձ��y�ձ��y�h4�h��*mu�)LΧh4�h��*�M�1<5X��[5:q�E���Q�!�`�(i3���q`�x!�`�(i3!�`�(i3!�`�(i3�q��@|�!�`�(i3<�6�Q=Ōw��QH!�`�(i3!�`�(i3~��c�'E���Q�!�`�(i3!�`�(i3!�`�(i3��]��;�nsȸ�"rR!�`�(i3!�`�(i3~��c�'��~ǳ�!�����(�I�?g�f�ja1�n�[�c�/�O��?�;��XC��o��y��9�ĒTC��0��$�>��w�����N%
��̥㡡�u���;�Թ!o�o,%H�%�p��� ~�/��_� H�C�I-�#��h`���r�O��C��0����bm���?������@�����c�J���<�"F�6x�_uS�CO�����U���o)��W�a������qθx���]8d�\�:H3?��n���N<�n�]��xw��猅
�V[α)j�o�R���V�8yd����Eg�~p!ۓN<E�����@���ަ��%�|%��]
�V[�圉��`�q�r¢w`�&qQ��00�c%���]>�x!����<u��w)�S���f��^@�~篟|�<8�F�-:��ԧN��78�:r&@��$�9��_,n׎ ��73��>g�����Mp᫼���hvK+�va��2鍔�	g\A���V�2���y�͌�4r�O��C��0���M�<lbtss߬����M�!�֓��u���;����\_�MX�9�I�[��On�AN�.5f$��F�Ŋ�����}�K{ɈC`N�z����le�kI��Ř�^~tҦ,��_!���5�NnZsA���r�O��C��0��D�[T�Q~�K��fC������S��u���;��l)P�u��F"lܵ^��UŚ�p-�q��F@�u��w)�S�3k:�(�-����Φ�AȨ�)���~ܾd���Hߵg�6�:���&~ZxV�3N��f Q~�=V"N�^{")8�*I��Ho��ݖ��u'�Ҁ��|}J���Z/��J]�j�j�P��se��^
c������Z��Ӻ������7�FWY8�{")8�*I���]^SΛXV奖ܕ��RL�a)�Vu~c!��,�%��WȺ�V��y!�M%��6�u���;��I�6r�����N�>A��@Q�BZ�n�qD���[U���zE��p��qx����-&���#��1��8�(�R/C((�%A��I��ך�6`���`i|�o�߫��<!�f�2m��u��w)�S�3k:�(�-7��Mv�9\��(
�m�ó(��8�:r&@����p�T�c&�׸P)o�KӜ�u��w)�S�5� �p9�AE�t�ݙ�����m�w���P"3��
f����jR�"�H�ٳ,�M(F�N��d�>�l;��r�O��C��0���/���k���_0��*�Ε�u���;��.~�Gj'��w9����`e�TS�?^
ر��ZXty���`�c�~e�0�We���ܮ�c:��1��q������-i����^!`w�� ��A�]�B=>_�o&�8��/M4#>Y��<<�٤:�e��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcUz����~2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��r�����A�F�7���3�GXS����E@��~���($�J.���
�=W�֯��i@F�5�=h�GD�#�̔"v��ƒ)?˳R����.��ѬL�1m��+Y#_WӢۉ���2=�l����ј2��<���,I\�Z˻r���V�>!�/�7��u���nEA��"0�qv+6�Pr"?D2BC��5��Yk"1/���%	v3�Dc�c~O���%H�$�DC.5j��?�y��hBQl-m
��	���q��q�©��'w��
�f��]�/V��X���V�2�Ct�z&��ÃlO ܅d^�R@Κ�2���ei"�,�>E����\�vňu�,�s�^�R@Κ�2�l~�Uf���}��\�v�T?�7G|`�UxHj,��|��	�"�,�>E����\�vňu�,�s���2��̪U��֜��3"�,�>E����\�vņ�Q�]�ޔiyV�[R�^Ƒ��!�`�(i3JHn��z�_c)���8���bg�1�Z���=�������b9����,����d���z���ߘ�)�I��<
DN�l0��F��j�q	k���A���������]c���H������i�=]A��O�T=�4e=��-f[� ��³��w�[��C��!�`�(i3���D	��U�l>o��|�,+$\�M��wF4��0[����	��N�Ae�#����ꀍ!�`�(i3c��Et��q���U����?�!�`�(i3Y%T��BPe.��xu	�>��l%i�-�|�)՜�4!�`�(i3v�ј�"��Z鎬����(��eظ�_--���g&e�l�����-��%Mm�jp=�>��o�
�v�ξ������ei]��fM?R�^Ƒ����"X��[��Q[R�7W����GS�*;q܄}͟PP��Z鎬����
C��8q��f�kN�ı&l����G<�e��
T�v��1���6��	���`y����ꢤ�OgZ)[���F�����E��@IE�U��n�-�6��
�jW��D���M���R'),��`��{|*�"��i�_:���5�%]���a(􆿳�ؖ��d�I�� �:&��I�?g�f�ja1�n�[�c�/�O��?�;��XC �Bʕj0����67�a��c���}��D���(��z�j�)�q��1�:�Ω�=A���>�LZ*IV���^�������m�q�,⏇���;�z*���Be�2l��4�y��ɦ�@^7&ģM�'n�^0o�<:�W�_ĵn(���˧�0z�cULjaGkƊ~F˯�+)�"j���b7|#9���hY����r�{p7�j�pܔp�l
d�o�R�GI$��ǂcY�~�s<��MR�������c�A�L'G~��6�7�5�%]���a(􆿳��?ƾ������ ���U�e�7����	N^�U��J��"ї>п�p=	�˳͠m�xW��9u$d9�cx�S�����S8�����NlU����z~��6��	���`y����@����gG<D�n:3M �[e�~'��Vh���*ܑe�W����n�4�{lGD�V�B��иܖ��A�.u�r���,DTc�~y��i�i��욕�'�e��`�)�	�%{�;����f�kN�ı&l����[}�@��L}�
�?�$���]׽�"�,�>E��0!S�,��ш�A3�(N��㎏qló�@qS�����8��';�¬pX�徯8�2�J���!}�<pI�*P�?��{	e'2��p�m~|��8yL2�����ތ�1�"5� �S�n���&&�F˯�+)�Pg�����R�^Ƒ���P4ǲ �n�/?S�+���LQ�Y��]��I#^�������8��'��������g�,P�n�BL�Jx��������k�V�6IWJE�$��dg0J/��=��K�E��{#6�aw�"�HߢI|{�0Lʡ;�¬pX��g��U-�ez�r�6��DP֞ �����Ə�_���ބ6WpH7���
I@1�ؠ&���Z02��`�z��GZ>.�0�i�ܰAb!��u�mj�B��V�}0�z��[��Q�՝�i�(�S��]Q�I����踫g(�r� k�|6�8-+��B�G�
�CӞD��]�)g��E����F�BL�Jx���`t�A~�9�{u�:�髊}���ۋ.�?��u�htGW�PA�;�֋`N&l�����*����s��'>s�a�x��{�6�e���ӯIJ ��`y�����g�,P�n����|!���^��\i�@^7&ģM��i;'~��% &gp�	8���R}�
�?���R��M�e.��i�X�_�0��'nUQ$n�ti���#M&�4�q�Xx�=�r�e��\
Z鎬�������(��<+���U�"5� �S�֯.I�ұS�)37J*uc�A�L'k"�jСN}�m��{B���T�D�]�!��	Ǹ�y85��ZlG���g��U-�e�{g�w-iI9�o����"��y= +i�1�[��Ka?Q�lXw�X�*xlL��I+=5�zߴ�� h�ҩ·��L2�nק��ׇ��r�A$�_�n��[��K�=T�_mQ�ǌ nqҺ�Ie�<����="�����:��HN��R��bP�63Z�t�U���G��&��/Q�g��U-�ex����焒��Հ��P���p�=̓�0�E��Zf[� ���-����5�����}Y�]��h@�Y�<���Ŝ���>�3I!l���	�|���/��@���#��M&sǚv�j�����{]F"���%>�rG40�RS���$
�)������SENan&��Ąk��msb�d"L���uL-���N���kb�r!�`�(i3�zk���)P<�ܓ�Yfĉ>99��R�Q���~�[�޶�r�ppE�"f�;�P�t�5�37y������(�;-O�{��&�EE�ޱ� p-�a &r|z݃3��윞+�5 �>��\p~z�r,$
p�a���Z��PlJ�M�=�혅vº�w�⽒���M��ҹf�f3';��|B���r����R(ǜ`���IX0F�MV�ҁGG�.Mm-;�!�`�(i3��èV!�`�(i3�'ž1�|�'����u��r��!�`�(i3�<��>��h�EtC�<�b_X�XV�b�z'hۉ)��d�7�q�!�`�(i3W����GS�*;q��=<�6>e��0�U+�qbp@�!�`�(i3`���*1
�:qEptiND�S���/9�=eSe.��a��o��ѵ��.�~<�Ɵe�*|�÷�Wе !�`�(i3�s�Yls��8��GM��-����!�`�(i3q�\E��0�����?uA|�d��?KYC'v�}M�9s��!�`�(i3��.J7h��r��H҆�.A`��x������D�f�6l�}��}Dq�f����%>�rGO�D mWN!�`�(i3�5ߧE4��!�`�(i3��ܐ�}ħ@�BY����;b�-�2�V��	��y>�����HN��R��?�d���&��g�]Wt~��^�V!��� JO��"�5��Dz�͒�p��e"5�O�%E#Pq�\E��0�����?Fe��1������Ə��}Dq�f�mj�B��V�-vR�Ψ������S,��!�.�g3ZE��g�Hb �;�����=��YV�v�\�b͐�	}�@�w��˪?�-���ei�^�̷ؠJ��:�����U��c̫IX0F�MV�ҁGG�.Mm-;�C>��ӚH�RtV�^�'ž1�|�'����u��r��FwZNE��=<�6>e��0�U+�qbp@�՝� s�#04~B3��������h��`�����y_�mS8<�n���F�P�7��S��h��d\�����l��=�O�-v�*_�mS8<�nׇӭ���H�����0�و�@Q�kj� �v�қp ���C�ˤk!�`�(i3��4-劽51�X�c�rs�i��]S���D�'�)�Բc>ݣK�6<o�)�/����O��]��MԵ�x3���ʗ�%oc�����!�`�(i3�Y8�J���sȸ�"rR-��ټs�  ����'Z鎬�������(����.��$��Rfł��kS�*;q�ց������b�Bϱ�mj�B��Vh�EtC�<��R@��"�!�`�(i3���F��O��ݚ�Н��/�cLb���/��C[��'�)�Բc>ݣK�6<o�)�/����O��]��MԵ�x3���ʗ�%&vY��;�fĉ>99��A0ok��$f��_Ub��7��G_��$�)�vx��������;_��8W�w��fD2�es~�cb�P��혅vº�w�⽒��8�>r&��H�ʱˡaf)��;��|B<&ǒ8�|s�g*n{��`�e�%R�4���ة�~�y�w�.Y�[���c$��oȺf��j$0ʽz�a?�d���&��@��v{�G[�8Ro9P�Ʒh7ܟˇ^�6� k�|6�8��tl2w�e�W+��W�FkH��۟�z��n�*�&�v������⪂!t-�u	D�&��9o�d�E�"�m���rwӷ9J�E[�l��a+Ĳ
�),�#�T��6�"�m���r!|�α+SƏw0��C�ݥc&�̢���>�W��*(��3H��ieLb)�5�o�' ���@�0�0c��L>�W��*(��3H��ieL���]Cr$' ���@�$� %7䨉��%>�rG6j�"Hsʆ
q�8"�@��v{�G�U��k":�ct�0��3��O	�T/ k�|6�8�a"�/A$���Z��!�`�(i3U�~�vmȋ���OH��c���鿋�E~��k}����/C.�L:,�s L�Zl�W��{��]�L���/=9'�����mC.�L:,��i���A��ݚ�Н���hY-N�g3�)��c�{I���,'�*;���#�b�>{Z����6��.��Lj�)6)-
�.�g3ZQ�ͼ���݌0 ���hT*.�Q��	�.8��5X���иܖ����S�f>x�:	�W+��W�FkH��۟�z��n�*�&�v������⪂!t-�u	D�&��9o�d�E�"�m���rwӷ9J�E[�l��a+Ĳ
�),�#�T��6�"�m���r!|�α+SƏw0��C�ݥc&�̢����{_8�Y��=�}�Vݨ��}Dq�f�����,�ǰE��C$��C�Y�\�P�p��jN˭�ޱB0w����u���ei�j���s��d���!i��'T���+`��W#s�'�yq������<N߼�K�iN��VW!��' ���@�$� %7�!�`�(i3U�~�vmȋ��OY'�E�g�������(ӈ���m�r����I��)���W�w��fD��Ӯ�n�w�R���y�sL]~ц�]$�x��e��U¿k�B^�(�8{���@^�4���zȯ�;�:���W+��W�[�ɝ������+V$}8�W�.��A$�P������5d�Q'݀�=��`���φ��<�6�_��(�Vgs��%H���ݚ�Н��r$ɓǃl[�Ƶ�1tSjv���'T���+`��W#s�'�yq���nF���<�W�.�P�	��
�Q�}Zt%��m&<�P8��PS~B;�T�dN�<@Iv��nt=:��:5A��p�̢k���F�KD�Vr[/}>5��0�B� �b��!�`�(i3y�}�6f&rG��Hb� h�ҩΪ���l�� ��H3�յXg:�$N��GZ>.�0~�{ ���ݚ�Н���'T���+`��W#s�'�yq������<N߼�K�iN��VW!��' ���@�0�0c��L>�W��*(��3H��ieL�X+�' ���@�$� %7�!�`�(i3Zt%��m&<�P8��PS~B;�T��Q׭n�L���/=9��9����C.�L:,�s L�Zl�W��{��]�L���/=9��<��&C.�L:,��i���A��ݚ�Н��Ra])n#�������k#���&l����$�<�F�q��-����!�`�(i3FkH��۟�z��n�*�&�v������⪂!t-�u	D�&��9o�d�E�"�m���rwӷ9J�E[�l��a+Ĳ
�),�#�T��6�"�m���r!|�α+!�`�(i3!q��V���<	s/.�Ss�g��+˘\5���jmY�VS���g�n�{�6�em�;���!�`�(i3�k��^�1gO .��0w����u���ei�@�ܫ՞�� h�ҩ�!�`�(i3��hY-N�g(�����+�F�$-��,'�*;���#�b�PSK=�>���@]vK��L�'`N߼�K�iN�� ��t΀�+I@L>���@]��}Dq�f�!�`�(i3U�~�vmȋ��OY'�E�g�������(ӈ���m�r����!�`�(i3��jVѭ@!�`�(i3FkH��۟�z��n�*�&�v������⪂!t-�u	D�&��9o�d�E�"�m���r!|�α+!�`�(i3!q��V���<	s/����AIe��0�U+�qbp@�!�`�(i3HN��R��bP�63Z�t���%>�rGO�D mWN���%>�rGO�D mWNHN��R���IX0F�M���`3�J�l��0(v}�	76�&�;��|B�6�'Z����Ct�g��^l�������A$�P������5d�`UNP�{y����:�*" �`�r$ɓǃl[�Ƶ�1tSjv�SƏw0���ĵ�%b_X�XV�b�z'hۉ)��d�7�qĹ߆�p�hؽ!�M��9�a>*<UB3 �~k�%����ZAL�:.�
9� ���(ٗ.;���JTv���H�����Yu�������&G!�`�(i3��hY-N�g,f�4w�E
��hY-N�gj����GU�~�vmȋ��OY'���}Dq�f���Ě�����}Dq�f��5ߧE4��HN��R���IX0F�M��'�v�|��;_��8W�w��fD�69|+)9x�����#��i7N�_�z*K��Q��O�بeD�I�E�����+T5�O�%E#P���_���ꪍ����:Y�{'%s	Hu�L	��E���v��&l�p�q,!����,�ǰ� Ϳ�&�vk	��+�� n`Ip�\{ف(�7���<��Y�&l������8y�Ɋ����Z���F%�X�ԼQ�}�p�?7P���`$�P.eE������v�h�g��U-�e a⣃_B7�}�!��?KYC'v1��E:z�'�=;v�����Ə*J�X�$��c��GlhŦ�.�g3ZrZ�0m�\�S��u���F%�X��/����7Fk����PqZ�o���ia������v�h�g��U-�e a⣃_B7�}�!���u��g��L1��E:z�'�ĩk(�CQ�r��H�*J�X�$��b���9C�.�g3ZrZ�0m�\�H�z��.�g3ZE��g�Hb麭�H�κ'��G3#uV��rU�w�⽒��8�>r&��H�ʱˡaf)��;��|B
y�3~;�>g��4� �㎿���o��D[�h��4o�ݪ����Vo[���˚����Z���2��}���/�^��;N�09h\�`��wd�F+��I��)���W�w��fD�?��+�|aT��3G?�d���&�'��G3#u���(�'�|�7����c