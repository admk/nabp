��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-K�趹���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�=A���>�L'jf-�6U�P�H�q}^���������g�3�7x��������&�ǝ�+zA��]��~ا@H;�W ��W�5�k��O��ڴ���WЋ��I�?g�f�ja1�n�[�ެT�Z¤��I^��?�;��XC��o��y��b1Ø^���#K���lӧIA�a�V��R�5K�yQb�I��68�/�YJ�'�دv)h�V~�$v�p��"}�vo7k2a��pP.S��*����طǪ�`DY��YH\��!���1R�_ߥ�]��4�:j�l�,9��)'��e�Ni�H�f���Zߧl4���0�?�1~�x�c�	�L}���i�m���w�*��O0�To��q
�-Hϭ�b#Ӡe��?�F��&��q�©��'w��
�fʖG�œ����s��3�mufҷGپ_7\F���r��RL�a)	�n-�~F\Y>;�>[��'�?�9�����9����E�u���H�nB0AܿҚ}�?��,9����	�ŀ�<J�Rz�5�Y�w����1*��w���r� ��<�3hY��RL�a)+{(y]&½�������$MAF�婨{X��ֹY���8]$�_4 ���L�A�k�8���҆�|n���6��.7��� 86!5��#�f�+���C����
4�
��|ſ����m����qB/������K0�m�!=�y����h�}��b�Z��������-?��1m��d��U�)�KD٨�2�&*����"E&��� �
�V[΋�L:�!#R�hgrH��~����й�I�ڔ������
B�u~SK���B+��b��?K�3�5Ὲ正�3@Ѐ���`�����f%%ep�t����%P�2�>�*���*��O�to���sp%II�~�>��RL�a)�G{�<��������O��w��)����cl�ֹY���8f-�.�f�*~�.��4Xy�Q��J�J%H��	m�Q� IA�sDqPGD@s�i�W�r����/��Y�{�ڌ�2�L�*6�	�\	%[h)�u��w)�S�3k:�(�-\Y>;�>���(i+�@1 ]\��Ny9����E��ű��k��'��^<?�V���#��X�*�& ���m:��@���i�d�~[�p�#��"SӠ�|&��yY�ao�;�z&�aD��/ ��è�ѵ�Th�f�7��t^��RL�a)ѻtUWR�������ǹ�5���L+ɓ���ZֹY���8Y�G%�H*7�"Acp�J����ID/��i*F�%�=����Yp����c�J�4�*�=�s��x-0����J������%���(4��AYp��t�jPP�
� �AH�}��� ��8���X4�c�$!sV���Hky*��kS�O1��l�t����@˾�����kx����̬���_����	x]́��D�^����i�6��87s�!��`�U�9�4 ��W�&�k�8���҆�|n����0ӵ�����ڒ�3u|?�J�Й�m�K�ţoAE�'E���fFcņB$�~�T�2�bT]�܊KMb�w0�k�8���҆�|n��1���N�N�SV [?/�����W o?�M��;]�#>fS�H��K��l��fu�Z��"R��Hv�|{")8�*I��_YLw@�H����>8��\�����^gF���0r	+2MWm�Q� ���,�Nk��6S�䥭*����	�z�}ݢ�Qy�?3�Vǡ9���<aDK�^�aum�Q� �8=��,�}����;�P���Ħq�e�����4�})���\�4�sg�oXx��U��������"^Y怄FUR�.�;�~�MUs a"�x���2@�+���c�#s�0���!Z:���:r�a�u�����!�M��E��ǮZ�`/��aG�k�8���҆�|n��/7� GD�����G��F��=��J�Й�m����ǥ�P+<�F�z'�_��z�Ӧ�'�b+aQ�wT�	$~j�u?a'���]����Ϭ	N*�b��n.�G�@���y{��O2��@����ا�k�8���҆�|n��]W Z;��T�ƚ��Թ	SL!�C�J�Й�m��/K5r��!����%�������Q���K�u��\�4�s��u�@��)����+��JHf&k;�F��o?�M��;]�NT[T<c�r��b�q,S}�E8yd����Eg�~p!ۓ�."#�$�.�x�Q�\g����>�`+ZP;7��
�+�0�6��z��ԊV��G� l���Q�r��yû��]��0gg�~p!ۓ�o�^�+}�D��"�Y�
� �AH���CdZ�G��vJ�^�Ry~�ҩ��N�]�J�Й�m�a�|goS3�K&�. ���Rk��4����蓻�?IkT˱ �T�٥��T�Sҥ��|E�EYZ/��>�&��c3�S��3ZT�{�y%��&��j��n�\�ys�}$+c$��笈������\�4�sP	�b\qB8Y�&�\�c��7�	eIW	I��?G�~�MUs ��z�~�q�'������[�m�~{��\�4�s�q�=Q��x
�ԟ�drȂ�~��]�s�h6q3o?�M��;]\V�A}��}���V���8e3Z}�ax�� 5�k�8���҆�|n���:�o�E��Uu-M�rt�d{��}lJ�Й�m��?�Vޱ������{����VjrHS�w�MH��j���r���+W��YJt�,�y"r� J&g~���c*& z�s�ђ�B�~f��0(�/��$ }2����T���Q���!i��ӯ�02�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vce��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�׍E�+��
���*,f$�7Q0- ��Ck�fÜ�2/���}����сsU%���n��/���Û�E�tw:g+��T��d^��_|��3g�ݜ��s8[Z�`
5��*�z�������D���J7"�x$�^w��ѬL�1m��+Y#_WӇ�s8[ZΑ� �}E+��)��6�$`=&��g���?��J��(����5�2���[@%����nEA��"0�qv+��r����N{a�9O��Yk"1/р�{:��'��팣+����F�N~Y�pXTN�v��ea�;y� ����t����M����3��~ �Q�^�y�zL͊�q��UG�s�����M����V�܄WD��|�����u*K6HT�����N�t�&_���9�!�`�(i3l0��F��j�q	k���Aj޽���Ǜ�����������i�l0��F��jT�����N�~ `�T�v��1��B�wj$g%Ah�%4
>��XP��Ȩ�wl��h�d�uY�؃�]n�� ���3�ҺIÙ=�H��ˡ�VkLs��dJR�^Ƒ���Q�^�y�zL͊�q��Yy�u'�7�;�r��0I� X�1��E����F���8�TP�}{�Z
M{2jR�j���m l�o�����зq8�Ј)w�<�_N �VL�(\��'&S�39؍��R��j�.(Wx*��|��pe���b������5	���]���>����C�h�'f R!�`�(i3��|g�Y�'���Xw�E�i�m}6�B�r���E����F��j��\w��0]EOJ�uxm�3���w�@V�"�����/�]�!��M8���	D%��_�ͅ��/��=��K�q�?l�_��ct�:��RE��W��_�ړ8���/��^����r��H�+k&v�Iz��j���'b�t	�U���C��O]r�<Uee�,�Aٺ�H�NI�:7�N�5�%]���a(􆿳����)T������ݤ�v�ϭl�\ѵ�Th�fܯ�ko��o�����}�ꢤ�OgZ)[���F�����E��@IE�U����S8�����NlU����z~��6��	�\�HP@�a���н�!	ozqP�"B��$I��w��,�������ݹ�0�������Dɵ�p�AJ�e�$��\�*P���8��';�¬pX��g��U-�eaԗ5��C�6�ǌ�lA�1�:�Ω�=A���>�L'jf-�6U�P�H�q}^������kK�N��ī��r��X/��4�q�:�"��yȯS���Qߵs<��7�m��+��jTʱ�:W���	�)�0�lOq��"R-��by��L���s�h�
!7<���������	N^�U��J��"ї>п�p=	�˳͠m�xW��9u$d9�cx�S�����S8�/ #O�)R�^Ƒ����"X��[��Q[R�7��z�h��4f��Ԝ�]����n�4�c_����+#��.X���*"v%)��Qcm h�]�!��	Ǹ�y85����J�f;�¬pX��g��U-�eAJ5ߝ������n9읣_--���g�vh�1�WpH7���
I@1�ؠ&���Z02��`�z��GZ>.�0�i�ܰAb!��u�mj�B��Vhs5e�U�Ͱ��Le�2l��4��a��se�ξ������ei^�7��u"@��8�5x�|����1�Z���=��of�-CD֧�ǌo�9ct�:��RE��W� y�T�v��1���2���I��'��{�6�e+Yi=��o�IÙ=�HVkLs��dJR�^Ƒ��V���"�VAM��n\�֥��ع���^[_�e��IÙ=�H��M����V�܄WD��|�����g֋�&l����R���o����$�1�=z�>���@�<[n^/��u�h踫g(�r� k�|6�8����^��L�de��y]/�qF��6��	���`y���h}Nw���U�m#j[3���w�@V�/�˟��7<���������	N^�U{xN��i>r�<Uee�,�Aٺ�H�L� s�j8��L���N@�/�M�9���{p7�j�pܔp�l
d�R�.��On��M��ҹf�f3'i3�|)sՀ�/V����!�`�(i3���^��=z�>����ep�G;w���w��l��ML�f���|����OxtX+�Y�G��"j:}��M�+����ei�}�"Io?�?��A�^kAO��t�+���LQ���"X��[��Q[R�7��iM��*����6*�Gc_����+�˂߮<u�4�!>I�W��^�����f��|�F7�_���}���.q��+����eǎd .8��K�Q��8��⢙���$��O�&��Î+,�C�ό� �������go�����h}����g�(tPw�uЅ�^̽1�� k�|6�8d��)V,��G&Tf��9x��p��;mQ��8���/�a'�<� \�� |+vܽ?�w-�e.��i�Xⰸ�7�K��0�mO)�}�
�?��(R\֎u�ZWž�C��q���U��@����gG������G�l.T��=ȵ�ixUS�`$�P.eE���lC��U�T�\ ���|.�Tӏr��꘳Uj{���*O�=�ͦ��]�C�K��ƃ
ᾆ�x�T�\ ��i3�|)sՀ4$`8aq�W�� ��uSP n��"����1���5�%]���a(􆿳���2����.ҹ���+F�]�5LdW�Q�����9w�gs �\1�Z���=�"j���b7�������B�D�F �ƥ�졪�Z.��0�W'���Xw�j�7���{�6�eυ���K���`y���pzl��a���JQ���8��.����Z鎬�������(�����9x��p�5��/��8���/�a'�<� \�� |+vܽ@ E�����d�٣��c�A�L'�ٙŧ�)#'6���;8=�g��U-�e�ˍ[L/}�t%>^�ߒ.�qO���WS���
��ٴ����9K� 	�c��#�6����]b!��u�^��po���s��d�\[]Ǒ�J�)�xVR�Hؑ悍!��2J��`�ѐ�{�_P]��.e���2J��`�љ����\������?XW�~a���@=������yM�˴�p�A�?�9�e�Dcb��܏� �� +@��睅H�/zP���o�8"��nH9�ئR'cf���a�	& ��?�d���&�Je��0��-&�6��_���9�����d�J��:����(Y��:���R'cf���³5��&l�����#W�U��ظ�d���!i�/��@��C�G����]'\gWg��	�Z�kfc��2���8[�����(����<m�H����Qw�c4~Nr_�mS8<�n�ݚ�Н�?V��j�c>ݣK�6<o�k��G<Y�dN�<@Iv��nt=:��:5A��p�B�'��a� 7�J�[|�m�ߕ�E�g�������(ӈ���m�r����!�`�(i3�k��M��߆�p�hؽ!�M��9�a>*<UB3 �~k�%����ZAL�:.�
9� ���(ٗ.;���JTv��!�`�(i3y�}�6f&rG��Hb� h�ҩ�!�`�(i3?KYC'v���ʗ�%���S�*(�����Ə!�w(�y?!�`�(i3��nސ��3���w�@V�  ����'mj�B��V3�����n!�`�(i3$f��_Ub�F�S�1 �fĉ>99��A0ok��fĉ>99��φ��<�6���%5)RHN��R��?�d���&����yϔUw�R���y���,!��%.gW>�a�ut�0o��F�5(��~�q��a+��bc�n7�}�!��?KYC'v���NE!/ ,��rQ�i=�d�ЈH����@�/�M�=t�z 7�J�[4���0���V��	��y&Qe�}�!}�5�^AI6j�"Hs0vZ��ҹ��g]�)]+Ý�~��:���HՋ���)~a���@=�y�z�����?XW�~a���@=�y�z��U���!=UgR� �ұ+s�Di�R{{���5�&_��s�֙�-���^D�V�{�S�*;q�v{��lw	�,Bp��S�i`YS��� 7�J�[���R��u��g��L�Ѧ���w3I��P`�k-:S�4��Y�Y8��t$��ɒ
���K�֞�`,9�H�W��<��Y�&l������8y�Ɋ����Z��t~�H
�)Ú�'nB�Qטg�u2Y��Pv����ʗ�%���6�7gE�s@�@�/�M��C�x��̬���	p�U��c̫IX0F�MV�ҁGG�.Mm-;��c�n��Xյ[+8�po守�ubs��2[�a��o���H�RtV�^@���~$�  ����'K7͍��|��W&":ȓM�Me���`6X��Aj��t�35L��$
8��2�ֈe�cN�0��ž�Ć�T���7X���c�}��po守�u�,l����M?��y��5�Q�d����l��1bx�cF�����Of[� ��2�]�<�k��u��V�Ո��Ú�'nB��!���c�A�L'0#P�O�Rfł��kS�*;q��
�7Cv��L�*dgN;�r��H�?X���V4&�zʖ>��;!�`�(i3�Y8�J����B�I��!�`�(i3=��,���H̷_��yC��S8�\�w�4�'�)�Բc>ݣK�6<o�)�/���C�$�ߜZ�`.��53���w�@V[Z��.�~�5�Q�d
�:qEp�;�P�t�5!�`�(i3���D�&��&tS�D�]v1�_ُ�����Ə?X���V4&�]Pn��J�:�_q�pWS�*;q�&l�p�q,!<�6�Q=���F��O�ȓM�Me��&[�x�R�"�,bxqX��׹��7��~���-՝-xC�;��|B#���rM���p�8����~��VX�P��/4�O�V2y/� LB�}A�
�V[��~B	G&].}&(�������\���b�dh��η�
��v\��� ck��`,9�H�W��<��Y�Ǚ#Y\��?�l~�U���� G�_��s�֙�wvA�qS�F_���ٱ'W�w��fDfTYQ0b| ��%UG�f���ՆBq��!��Q�R���F�(|��8����ei_��s�֙7�}�!��!q��V���'�Pp��XO)�Q>�W��*(��3H��ieL���1��#��{�6�e
��>�i�g��+˘\5���jmY����A�I�{�6�em�;���Zt%��m&<XdYʼل��OY'���c���鿋�E~��k}����/]P�����+���LQ����$�����E~��k}����/����g�p�+���LQ��:5A��pw�R���y��[�ڰ��7f�ڭě�m������G�
Rv�@/�uw)"/��=��K�R��K<_8 _��s�֙7�}�!��!q��V���'�Pp��XO)�Q>�W��*(��3H��ieL���1��#��{�6�e
��>�i�g��+˘\5���jmY����A�I�{�6�em�;���Zt%��m&<XdYʼل��OY'���c���鿋�E~��k}����/]P�����+���LQ����$�����E~����t�������s!��"�m���r!|�α+I��)���W�w��fD��g<%���]c�T�Ŧҹ"��s�D����_ �Q��ǺΕod'ٙ� �z�:Y���J��:����SƏw0��N�ijR'�yq������<N߼�K�iN��VW!��' ���@�0�0c��L>�W��*(��3H��ieL�X+�' ���@�$� %7�!�`�(i3��`!�r7q����1>� {�}���my$�N��o�/���;fĉ>99��;��|B3���Hρ��~�_�=%䟳��L� *NK��阬иܖ����S�f>x�:	�W+��W�FkH���8ч�����Dn��i�Q׭n�L���/=9j���)��Q��\@
����G3҇
��'T���+���J�N�#3�)��b_X�XV�b�z'hۉ)��d�7�q�HN��R��?�d���&�Ɲ{�N� ��Q:�TO	�~����Q�y�$��A$�P������5d�`UNP���èV\���F�`yx�>�+X�M?��y�!�`�(i3��8���L��Z�|E�g�������(ӈ��Z��&61�7���'S/��%D`����AIe��0�U+�qbp@�՝� s�#04~B3��������h��`�����y_�mS8<�n&���S�RRǚ��ظ
��@�U#;�jmT�#�,l����M?��y�!�`�(i3����o�al&����Ŋ5�m�XdYʼل
4�e �S�{�ܦ��ܶ�iD.l^S2t�N�/�ڣ6��:[+b��'�Pp��2�!�,�
�:qEp�;�P�t�5fĉ>99��A0ok�׹�� �ѕC?"	�~������*j p�⫎�`ru���L}�sL]~ц�]$�x��eC#/<���q^����+���@/�*<!�F��66����~�fE%*)�匥��m l�o66����~ω(�$V�y�2�x�h������M�!��^��BcƬ^�)pE��d���!i�� л����`3�Jg'X�~bw��U��)���Y;e�iK!���d.�� л�{y����i�q,?5q&kT҉­���+V$}8�7�I0I/RR���Xc�Qw�c4~Nr_�mS8<�n�ݚ�Н��B�.�4Ӭ�P8��PS~�Dn��idN�<@Iv��nt=:��:5A��p�� л�U�~�vmȋ��OY'�E�g�������(ӈ���m�r����� л�����g�Z��3��a���!@�f")u��r��<�6�Q=y�}�6f&rG��Hb� h�ҩβ��y��lD�����U��.��r
���иܖ����g���u��r��!�`�(i3Z��}	���C�ݥc&���XO)�Q>�W��*(��3H��ieL���1��#��{�6�e
��>�i�g��+˘\5���jmY����A�I�{�6�em�;���!�`�(i3����j��`��W#s�2t�N�/�ڃ����<N߼�K�iN�� ��Tv-_�0!>���@]vK��L�'`N߼�K�iN�� �Ե�����,>���@]��}Dq�f�<�6�Q=��i��:q�M� Ѯ&U��8�>r&��U�����Q-s�H�RtV�^!�`�(i3�ٻY84����<	s/S�����g��+˘\5���jmY�wΦs� ��6��.��L�la�F�wF�,'�*;���#�b��{�.�t#6��.��Lj�)6)-
!�`�(i3Z��}	���C�ݥc&�̢���>�W��*(��3H��ieLb)�5�o�' ���@�$� %7�!�`�(i3��\ NhA� ��_��5X���иܖ����Sp��;�{��!�`�(i3<�6�Q=��hY-N�g(�����+�F�$-��,'�*;���#�b�PSK=�>���@]vK��L�'`N߼�K�iN�� ��t΀�+I@L>���@]��}Dq�f�!�`�(i3�ٻY84����<	s/����AIe��0�U+�qbp@�!�`�(i3��\ Nh'{w#/ B!�`�(i3Z��}	���C�ݥc&���XO)�Q>�W��*(��3H��ieL���1��#��{�6�em�;���!�`�(i3����j��`��W#s�2t�N�/�ڂ�nF���<�W�.�P�	��
�Q�}!�`�(i3��&.��8�F�S�1 ��� л��5ߧE4��!�`�(i3��&.��8�F�S�1 �烉s)�v��IX0F�M���`3�J�l��0(vC#/<���q����,�ǰ�L}��tO��*�O�{��؉j����[�O6�o8:4�I���c�90�Ǘa��xO.C��WHe�Q\���F�`yx�>�+X�M?��y�!�`�(i3��8�Zⓞ��mdN�<@Iv��nt=:��:5A��p��$���͜P_�_S:g�RMm�o��'����Tj��^�G�E�BS�+��U�,�P!6���r����܌;���'����u��r��Zt%��m&<����Tif���G��8���L��Z�|u�L����'S/��%D`1�m+�D8fĉ>99��A0ok��$f��_Ub��7��G_��$�)�vx��.��v�]���B�Ŗ��!ѡ�ĵ�%�%��L�V)���y{0��(�������M�!�OY��4q
UǙ#Y\��?�l~�U]R�.3N1z,:[b?`"E&��� �GM5���6��Y��\k�\�a�/3;��|Bﻍt����-�����#�Y�Cφ��<�6�@a� ���N���������y��o��7�;�jmT�#bs��2[�a��o���H�RtV�^�#~.��,!,�:�� ���?R �K7͍��|��W&":�;b�-�2�tiND�S���/9�=eSe.��a��o��ѵ��.�~<�Ɵe�*|�÷�Wе !�`�(i3e<�Ia��la��o���H�RtV�^FkH����T����!�숫J��M-03�gM�¨ɢ~2�
?��,��*�B}��F��
�:qEp�;�P�t�5fĉ>99��A0ok�׹�� �ѕC?">}���� ����!�m1�H���W�w��fD��'m�Yz,;7��"U�ag�ˈ�	y��ы>�~j�x�`������.��4�F1���l혡�s�5��LS*��ud�H�V�܄WD��|�����5+*�Π��yGb���)�tm�&C�bz�h�����.��4�F1����jaս"�f>x�:	�#��'J()�I��64���팣+�����t�T��?E-h��$^(?��"��h��w���`����k��M��'ž1�|�'����u��r��FkH����T����!�숫J�dN�<@Iv��nt=:��:5A��p��$���͜P_�_S:g�RMm�o��'����Tj��^�G�E�BS�+��U�,�P!6���r����܌;���'����u��r��Zt%��m&<^{ʓ���8)���� �X?�Vt��@���.#=��n��팣+��!�w(�y?fĉ>99��A0ok��$f��_Ub��7��G_��$�)�vx��.��vذYC�8����g����<�c�����M�~�E,��B�A��RN�-#���zym����HG�e�#=ذ{	���h�U�p��ٰ�Ř�hF\F��y5�N��b�����C��iF63���ш|m�Q� �ʐ~����R�"+��z޳�����8�{%C-��SL��@O��*'����N�1r����P�R�Ӛ�2i�F ��%�^O���EID$3���A��S6�w�*uI�2E���c7�t�~�<ͯ�G��R'),��`�a"��-K8�[|Un֥��ع��������������Ʊ�_�eD�I�2>$�]�U^���\�}A� SY�O_'�
�y<xІ6�I=T��\�'�`�'�ؗ�ly���@X�}�-�a�)�?z��3�kt*^����ɰ�U����NJ�q)�c��D�C���,���Ъ���\�rҖ�A$�P������5d�`UNP�{y����:�*" �`�r$ɓǃl[�Ƶ�1tSjv�SƏw0��,��*�BG��8ao���'DV���b�z'hۉ)��R���v�ء�����6屍K7͍��|��W&":�;b�-�2�tiND�S���/9�=eSe.��a��o��ѵ��.�~<�Ɵe�*|�÷�Wе !�`�(i3e<�Ia��la��o���H�RtV�^FkH����T��������a��&k@C�Ɨ0z�cUL��Zi+�E�,��*�Bkr���P�b6��.��L�=��gr(Ƭ�:<��j{�ܦ��ܶM������)̷_��yC��S8����ڝ��t��@����Yմ�nJ�|m��g��U-�e1�S�����fĉ>99��A0ok��$f��_Ub��7��G_��$�)�vx��.��vذYC�8����g����<�*>�Ƣ��}K�����nc+��T��`	��
�+����/�!��-`����7VV�{pQ;�im��h/ŭ̪��W& s���X�PC!���k��$���X_pU��֜��3��t�Bf{��dv��oTN�o?`��M�L����\7���JQ���8�Q&2TB[�л���7�0ݸ�w����;;)U��N=�$�
~J�N,�#OOJd֯&��s���qz�Gb��P���|��p��PIQ#�C,0�?���D�wP�/�w,/���` ́�x���������'J�I�%��Y���#�����.��4�F1���Gb	l��c�����u�6�0��ݫ&�b%%7���c��;;��|BN+-����]��.�Z�eր��������='�����|u���;_��8W�w��fD�69|+)9x{���Ej{���*��c����	�����E����k��$a(􆿳�cof��7��ܼCI�_���a���$ϓ^{ʓ��!wZ����dN�<@Iv��nt=:�
')���#�^�
����c�Z�~����)z`Q�.)�:)f���`$�P.eE���lC��U�T�\ �͂UQ����Tx��
�0���U! t"���9a�Fc�����l�����5�%]���a(􆿳�cof��7��ܼCI�_�����!���["�l@>�%HƔD:(�֥��ع�����e,w&�#g�k��c%�X�C�����V��C��_K�H�%�oT���tU�bFPs_*�GqW�w��fDQ(1CU���Z���Z)[���F̷_��yC��S8����ڝ���T����Isŭf�ҿ�Ʊ�_�eD�I�������q���6�6����D5�|أͽgF"?�Q��ǺΕ�f�f3'_��s�֙R���Bk�d���H��H�2��z�b�4��Ǳ߁R�^Ƒ�өwo��Z��Ac<�p{�5�O�%E#Pq�\E��0����E�I~�*0�ŷc?KYC'v�����G eK�lݧ}�	76�&�;��|B4<d��
~�_��.��ϕ��q�"��Jl��q<uiF=�xo�R�^Ƒ�өwo��Z��Ac<�p{�5�O�%E#P�G�dE�h����E�IȪG:vmX��u��g��L�������<�^._�}�	76�&�;��|B4<d��
~�~���.�;��|B31F��~m�>[eb��/��RU��H��<�C�Ar��� ����Dɵ�p�AJ�e�$��8y�Ɋ����Z���|����J�yؕ�o!�'��x��M���U����z~5x|���MM
��,=?�d���&�ȓM�Me��j^��n�_.��45��LҺ_.E��p���V�֕ߝԀ�3I��P`�krZ�0m�\�w�|J��c�ˆ�A��6j�"Hs|��^�p!"���(�ek��m6[��-�b�+�