��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-K�趹���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVD�6�����;��sD���L�S5H�j.F����g�3�7x��������&�ǝ�+zA��]��~ا@H;�W �v#��s�8��yW��V�>!�/�7��u���nEA��o��y��b1Ø^���#K���lӧIA�a�V��R�5K�yQb�I��68�/�YJ�'�دv)h�V~�$v�p��"}�vo7k2a��pP.S��*����طǪ�`DY��YH\��!���1R�_ߥ�]��4�:j�l�,9��)'��e�Ni�H�f���Zߧl4���0�?�1~�x�c&	��/v��ȭ��J��n�l�� �j_G?�8�E�A ǢC���s�7nF��%�h�����J�26�kk�`Ŗ�M]!ۨ"�`8�|=1|Y������w+2^ݲ5_X�� B̄^��R�8���2ObUZ9�ٵu�����!�M��E�L'4�����6��H4�
� �AH���CdZ�G��vJ�^ <.���fR����J�mJ�Й�m����
|H?t�sa��S����#���<Ī.5Y�`e�TS��\�4�sP	�b\qBTT	q��$W�7�>�Ė���A�r�~�MUs `��'�� �jT!�K� w�;�d���N�tכ݁=9�|Z���ߐ'�[�Z���1VU���+L��h��X�vB#|y{����P7�.yt�gU*Z9B[�^������+�ͫUz����~2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcMD��y�sY2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��(M�vS��~�X�x��S|��}�ZC��aNvA�;�m�\��qi��p�7��Z鎬�����R�LM�e�IC�_�\H�F?t�)�Y¹w�.� -��E�I�?g�f�Jm*)�m��+���%	v3�Dc�c~Or���q P�^�&d�A|�1�:�Ω��
�/�r�ѬL�1m��+5z�P�_X�I�?g�f�L#����2=�l����ј2��<��L7���%U�"sj� �<{g�P�r�|AڹDc�c~O%]�-q_�bI��'�ct�:��RE���|�r�HzL͊�q���a�����$��Xo��I;��?��H�MPq6.JHn��z�_c)���82��m �A?p\匔'넹GZ>.�01#��Z�����XP���3�u����$��Xo�U)+N��'�̗����d����zL͊�q��UG�s����5����`K��"~6���aq��qa�*���zL͊�q��1�KB|1<\�5����`KJ�	�LÆ�Ǒh�~��JHn��z���o�K�7��k'�w�����Gl�N~)�jA( ����_�h3��{I���s iG/Y�P	dU�1m���E�Y��Yc�A�/����<.+6J!p�m~|���53eT��@��]�h��؅��FJ����HwL�X2��m �A?2����u�ݯ�����I����8�TP����������s	I2��m �A?p\匔'뺪��k!��T�E���JHn��z���G7��7��k'�w�饋����Αǜh��6���C	)�H���o��qo�:�Ȋ+���42�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h��n>�ϸ����������&���$S�ݪ��1#��Z�����XP�����w�K�	�<���BSG�p�P9 �W	́�p�m~|�ַ��6�����=�$�Э��n8���ٽ��j�Q%��{S'��p�m~|�ֻb�UPM�H�ɇM0M�/�s���'n�^0o����z�C�f���v�+ʢG&q^�`
�c��><�$���|�r�HzL͊�q����$J����m��oK��BvGޣkQ�A���ۖ�{3�u٠��2���O���|c_�m��ġ��,�ɿo|��g�?� Zh�R?�R��n���TaZ/2��m �A?g�{�]4�W/S��8(�E���Kt�+Yi=��o�IÙ=�HvA�î��zI��'�����7���{r��I`1R�Jʡ\��ԙ��'n�^0o_
-��[��������p\匔'��Y��)�?Z����JHn��z��S3W�K@EU1��?��H����e k�|6�8�8��A	qhbvk~�#xs]p�[Tnn�.ᬵy��Kߐ��~�.E&��u��}�|�݌�ˠЋ�l�T�I4��欱���j���Ln��S�W�o��/z/�@����#4�5����`K��fx'v�ao.\C�k>l\��y0�$i��k��L[���p�o,u<@���%�3�F�a�si՝ӟQ��ǺΕ�����a�g()��ikp���H���0H�YS�T��ġ��,_R,T_<�3+p��@n7��k'�w�]a��1qh_�n�To�[�C��-��JHn��z�Lqܳ<��J*�Rs�0䁛����$E,�J�|Rf�� ��iԹ�08p�m~|��el�8�Ղl��=5;R�ˊ	18[{{N���zL͊�q����6���p�m~|�֚?��]t��R�}vJ^�j��T����'n�^0o�ߤ���!
f�Nd+l�Yҽ֗�+�� �L�������D�zY�lN�����&���1!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3<�6�Q=GB���mQ*�7`����M�Z���	]���.�#�.ZVRѿUJ��\���^�W+`�x�oP��@t�&�e�5
�`#_G����q�41&q^�`
�c��><�$��;mQ��8���/�6	�4bp�y�]�h��=So�?D��PL��O6��W+`�x�oP��@t�&�e�5
�`#_G����q�41&q^�`
�c��><�$�X~��\��o����׋��`y���]���.�#�k�:A�	S�+���Ăc_����+.�	|ǔ�.Yz�Qcm h�a�x�ct�:��RE��;mQ��8���/�6	�4bp
	�7F���I@1���t$I+�V�6IWJE�YY���F;�I�e�,��[�9q�Y�{'%s��.|Z���I7��-5���ӯIJ ��`y�����(��u�
_g��c��f�ܗ��DX<�c>1K �:;k�+��b9������|L�K�)x�?{���x.�Knqx).L����<om��N�+#��I��'�������.��R�}vJ^�Ԝ�6NzL͊�q��]� ���_�hbvk~�#x�r���sVnQ�rV�:uj�p�(7��k'�w��%=��ބn���㬺0M�/�s���'n�^0o�'vX[��vW4��`��?B��ž�'�t_� �e�7��k'�w��%=��ބg��� ��"Ki0j@$��U� ���_�ĕ|G���
|�NwWk�R<�����\���^�W+`�x�oP��@t�&�e�5
�`#_G�쵄����T�=�;^�6#9���k��$a(􆿳����^����z�h��4f��Ԝ�]����n�4�c_����+.�	|ǔ�.Yz�Qcm h�]�!��	Ǹ�y85����J�f'6���;8=�g��U-�eI\�53�fM +�gf�����w]cH>��DN2���!~;��i�̥%�CvK���9u$d9�}�NOI�i��h��*���RU����I��'�����3my���pC�f"��O�9�@��UF��M�5W�;^~m#���WY���
�_���R�p(��oP��<���yZ�����C�W��.hΕ���iv,�v�����&Q��3�ց���=�b9������U.6��`�ю龤9>(�vgx�y�Zgl/��mu��(��u��5����`Kw¹��<d���	fdLn��S�W�כJϾ�i�I7��-59�}
�lx��]�ۋ�މyFB0�;+�<�Iyp�m~|�֚?��]t���~j�1#��Z�����XP���h�5,Wl�/�O'�=�� U��k-I�!A(�����=�C��	:����Ȳ��%R�xsD@@&`�`��z ���pC\��� @1ܭ���U��+�Xa�H(�˕-�:I�x�//(f�|��*ܑe�W����n�4�c_����+#��.X���*"v%)��Qcm h�]�!��	Ǹ�y85�����څ�ɡ��ls�u°������Г������G0$�� ��U�E�0�LK�W�����Bb�fH/Ե,Bud�aZ��xV-����dN�#V��gUs ��ޛ_�.��k���?N�6�e�:r�"~oB�*v-��U<4�>O�6�ูS�K���2 ��4�E�>�����*ܑe�W����n�4�e��}i�eDI��'��d�uY�؅��|�r�HzL͊�q�����-������ls�u-c5����>&�&i���>)8�ӓ����J~�,Q��E�ʬ�_A�������s���K�+��uKE�WJ�2��m �A?p\匔'������^[_�e��IÙ=�H��M���o�G�m�?60���d��jT�������=f^I��	+�jÐ���g��7��k'�w�(�b�|�5�U����z~+Yi=��o�IÙ=�HW����vcyi��TrdP-e��h�q�G��S7}��E���:���'c_�J�p�m~|�֚?��]t��H�ʱˡgb'e�W�'n�^0o�!F�;^/K��^̽1���C�M$�;5M��)�Pt�e'J��\|YX�<I@1���t$I+�V�6IWJE�r���秹�3I^�v�[�9q�Y�{'%s��.|Z�����8��''6���;8=�g��U-�e �0$
�6�7��k'�w��y��3g��y����Z�� P��\�v��\aьIR=A�;�֋`N���}J�|���|������F�QY���=�w�Ηե>���Q=z����9�r�)۬
#R��XI��'����0/�e��9�S���ތ�1��\�v�?M-��6(uU����z~���V]��y���KT��$E�2��m �A?�����zP�����1#��Z�����XP������0/�e��9�S��8�U]k�(���B����_T���a�aq��P���F;I6�$��Xo����BɊ�y4<��!I�Ki0j@$��U� ���_��6F��.N�DMY����U��t��ܣ^\t�*�00?�9�f�u:�]X��w�3Ɇ��C��ǟ�q
_0�>˜��1��٭�*Q�<���@)�t�d�f�rЄzɳ�B��,��C-2�^���ij�IROgn�t���c5�V��On�5����`K�jV�{+煒�|�r�HzL͊�q����֒�����6:	�<�&|L�P�i.l�;�����.>m[��[D-�H���o���&�t.�}]���.�#�9�j���BD���c�c_����+#��.X���*"v%)��Qcm h�]�!���<C����5����`KiW��
�!C� �u؅��FJ��gm?2�I��6�]���~`��ʿ�ϞzQ��n��;��sD���L�S5H�j.F�>�k� G��7��k'�w�D!�[�[�K&�P
K9�.6��%���4]�k�1 �O�o�U)\�fl9�yn��3Ĵ�W�a����ڧ.��Ha�솒�T!��\�x3��2�	�4��'2۶��]=����߈���j�3�W4 Xy�O���b��0w�mL(��ߠ�����4.`а�TV�^Br�hM+�a�w�����W\������M{�2���i"���I��'��x�����m������7w|s���0�$i��k��L[����D��^'�⺴�/$�gۆ�F	ȕT�0���o� y���Dx�IY�'�ׇӭ��!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3���gAq�ޢ
v�@PFN�ؿg��i��ġO�/��� ���%�ћ��E����ׇӭ��!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3��jy4��8(��(����`�u�7��� K�8��?C�Ft����f�����4���s:^�y-!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3���w[�P>�X��1�3Y�/\�>�HF(�GϠ"�(k��� )���>�n��u�l�7��k'�w����%iz	�d$^���N�*}*���4]�k�1 �O�oT[¥�*|�·V��J�s�ggr+>��~�����~%��I���K8���]�BQ��zo��!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3&��潹i��'��\&v���O�1{*�	���^<�_��!��y��s�ѧ��0���൧&�~!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3W�	��tj���s6��h��@}Ih�ܺ�](��&�5�k���s����?�/C���Fz�!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3�(]:�z��ɲድ��L���9c,Ѡ�)*T��l@{�"ED*���k��̔�?�AXv��؄aX܇5����`K��|>������R�t�5�e͉�Xk����0��D�<T�kx�����V�Y�D?���'BWG����B��h�񿮬H��q�l�.iA�$��Xo���h��ߡt�.s�_i�k8�p}K<
4J&)��I��0:�Tm�Ğ�3=�ؑ����"�A�:�`Q�v��؄aX܇5����`K��|>������ROt+�z��e͉�Xk����0��D�<T�kx�����V�Y�D?���'BWG����B��h�񿮬H��q�l�.iA�$��Xo���h��ߡt�.s�_i��lS��4J&)��I��0:�Tm�Ğ�3=�ؑ����"�A�:�`Q�v��؄aX܇5����`K��|>������R����q���e͉�Xk����0��D�<T�kx�����V�Y�D?���'BWG����B��h�񿮬H��q�l�.iA�$��Xo�k�Ԧhg��������fQp�PU1��Q���n��̒��b�|ݠS��2��ò�{�"�%�F��CƖ�m��ֿ�Sd���\�� �*ad��%�Kuژ�!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3��[P1��tiV���ݭXIԒ��w��C(��{�_�](�U��Y�pc	�P>7��=!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3)�NO�娲Lq���2E�،��h�R�+F��ۯn����T1bl�
\����wR !�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3B��I�����\��RT�88�ӎN�5	F;������t�'2۶��wc��du˷�����9�G_h(��ۀk_��l0�$i��k��L[����𲱧ϤM�6=�?�i���۫Ex���n�h깳&.ȳ6u\���]P(���5��!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3��&�T�zc��8k:�
M6��b�h��7 O��Dt�A�4�%5�����=�8X�˞�DG!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3��D`?�����[�G�;�B����96n,V,4c'Y�s��f��K�D��ׇӭ��!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3!�`�(i3Y�D?���'BWG����B��h�񿮬H��t��;Pм