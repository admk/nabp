��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-K�趹���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�s8�R�	�}�����`h�ag������T�/ L�� ������[���a�8%`��4�s�6�XAoeuxLZ�#8v��fT��ı��¥���hM�,=i�@x_\q�jB�Fg�Y씤`��p��>�B�㬊�N����t-�!CB-U���T���딣0&_���X0���2|	p��rw@	@us���\���Z�
ۍ���yq�`݊�|���"rG�
���}�\�.�DV	��dU�;�\����vg������W�aeYgA���z�Ś��
��H,7O���u\GAݐ_�!����P�>���_�xEt��0��}>�E�(��s?��n;�|-���g]��~����B���hD���� ��Sɣހ��g�R��b�^��\�����2�����d�h$�;��I���*�F��QF(sOw*��kSa�����35}jS�<��,}e�_71��Z��G@� �O;��Cٯut=���Z�y��ʲrM��n�`���S��w�\�)ܶ3���Q\�_q%�~�v	�+h:�俧��j��R)djx�2�F��Ă�78�T8�+4ԡFZ�t�������ge�qZ��Xz��$b�[��|��\�4�si�W���
�ԟ�d��|�~��Q���K΋o?�M��;]O��c�D�(�V���h��6�h��\���2��m�!=�y����h�}
�ԟ�di�uZ^`3���:r{Ko?�M��;]�=��)�I��)܅��c�.[K��m&����~�CxT�Z�A�^u��w)�S��X3���7��Mv�9�C�q����k85U��8�:r&@���:�J��""J7��Q�4IS88+`VU��/�����J�|(��jrHS�w�MH��j���r���+W��YJt�,�y"r� J&g~���c*& z�s�ђ�B�~f��0(�/��$ }2����T���Q���!i��ӯ�02�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vce��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�׍E�+��
���*,f$�7Q0- ��Ck�fÜ�2/���}������]�0�lK'���Xwʈ���m"p�ئS��.V&��B֥/~.)��3\�R�F*}�c}��uO�b�^��\�-`����m�q�,j[�YP����M�g����!�`�(i3�E����F��j��\w��0]瑲��Zr�zM#��m�"�,�>E����-��%M�:2QYeƈ״$(�>g���0�&�ͭ�h�O�0"�,�>E����-��%Mό���.ӏwbk�$���7Z��!�`�(i3c��Et��q���U���
��I�PM�'�ghR�P��|g�Y�'���Xwd�n]N�/��A����Q[R�7J���hB;��i|�l5R�E����F��j��\w��0](@X~�H:6����Z9"�,�>E����-��%Mό���.ӈ�=�$��zigzA=v)!�`�(i3c��Et��q���U�ЂDa��(%װ$��_�zM#��m������
L'���Xw�P���w��:
1����s�!`��z�]2�y�Z鎬�����	�7 �# �����2�w�����|�Ƹ��]�!��	Ǹ�y85�����F�>R�wX�Ձ��̰�!w���B}s�!`��z��(�
t�ژq���U��d�b�ʪ%��1!�`�(i3�����
L'���XwI<��f�E�#D�����Ә�N^tӱ1R�m��+�<4��ˌ�ň��h��<�..�4��w�(�E* �Bʕj0����67�a��c���y�H�$�TE�EYZ/���!`���� �yz��$6�D��L���_�L�Ȳ�V�溜��D�,�H�Dc�c~O����*�+w�7�G�6�!~�"�,�>E���]�!����-ዧ�[�����bp���Q0�!�`�(i3�d�٣���N N�S�	�:-!@xNm���d�0x�梧���]�!����w�Հ�(.V��������lz|���~{�Z鎬������_�,��LE-L [_1�f���зq8�Ј'���XwI�&�\�+1���}x*ؐӘ��b����/�:�3�TF
%$�����!���d!�O��1��2�.w[�%�!�`�(i3�i3<�f�D.`�Z���L5ӥ���98�
x�?�����tz|���~{�kѶ���� ۹;EtS<FۈJ��R�Ws�N"T8�zn6�u���Q0�lC��ۺ_~5�Ǫ��I�&�\�+1���}xe�4޸5b+�����50)�}�����T��.��W����"�,�>E��ۦ� ~�p�+�����50)�}�����T��.��W�������E���b!��u�PQ�>\Ճ�I��b-���q�[���QR�hǬ�&Q���5r���$:��8ڇ�ȓ�iӚ/��E/��Fv��a���7��Z�/�Nc�?&3�7-��ԡ6���9�̪=����\���S)��y��숕iK�D�b=?#�ˏk����0��G��e���������6~��2��,u��T�KKnfO����&{���x)�o/�1_����2�K��n@�Xy|�WA�$�����jd�	�!�`�(i3!�`�(i3��+p��qR�Ovc�[��l�,1B��CSk�_�#g� |y��$ŧ���`3���jO����&{���x)�o/�1_���_��.)<��O����&{�6�LbE���jVѭ@!�`�(i3!�`�(i3�%ؙ,{F�2�����w$�Q!9Z;<�O��gC����hj���hɝ(z�ZI~,|,���pq�vأ�U�[�m��U��)���Y;e�iK-pm!9�>��n4s1�U��B��-|k������������r$ɓǉ�.y�U=������&G�7���������U���g�'�^����x��7�֕iK�D�b=��p�:��D9��ɰ���|e"��)�δ��Iћ<���I����~u���NM���(@X~�H:������宦%��s��u"���ܹ߆�p�h��d��JXl'�T��~��Uг�|<����&��m���d��(�[�*0��d`��������x��7�֕iK�D�b=��p�:�S1�ӿ�Q�ЙMǿI?����[jMQ���0���g�����;q	�%��6�W���b�0��%t̓�@�8��"�7ό.R��x��� ��2�w����:��q��5ߧE4��Fr��j�|��۞ͤR*̮؂���@������X7