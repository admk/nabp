��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-K�趹���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω�[@�qR�� (� ��"fف������L'4�����6��H4ي��2_)��:B!�b�ؐ:�{T�{df�r�<�XD�* O�:����>�ፑ���ԛF��W��`��q�©��7��#!l'���h�W��!��CR�����g�3��N�w	*D���y&�f��+K��[y��ڂ�1aY���~a1k��1�/lt�3� P�;��1�-���f񻲗��~o��:���F�q�\���z��<�Y��{^(�Ś��
��H,7���ZXWL�sZ�	!w���� �bRw�����IL�+�{Dr[��=�K)�*�-�>�����Ádo�dN<djY���o���F���e����n�QX�v����<.���+��T���O'�lR(���«�������d�ufҷGپ_7\F���r��RL�a))�kc�߇2S[�����mBQ��JZ��	g�_�Щ7C��H �!�fLfƇ������'ª�5�L���x�%��)􎺙�ޮ �-j$S�k�8���҆�|n����+��`!�"n��v���uWTJ�Й�m�BM�Ɋ�p��"�U��b!��u�>o·,��8D"�s�z:�Ebzi`Ht����	x]�fX�eϝ(�V��
:/,-���	�Ȃ�B�3ʦU�4C$#;W���]w t��������SۣF߱�y�Zk���GT�U�{�OJ%
������7%OU�z�z.��e���L�Y&Q�\7�	��,�;���<)䟓�~������ЎG2`j��Um�!=�y����h�}�_nR�� ޼pk�
�r�N�N��o?�M��;]�=��)�I��)܅�������1<���`z�X�a�������RL�a)ѻtUWR�N	:.���n:�ƨ�Ob�ky��Ǡ�7C��H-(�w�N���A����&\�/�� �R�+M��m}os֮7�"P3��_� H�C�I-�#��h`���r�O��C��0���df�� 0��]�������yW�u���;���A��j`��'�����`U+n%K)��k��Ǣ���N�y�Yc���;��sD���L�S5H�j.F�]^�t�e�{��/Ƽ���\�4�sW c`k�󯚚����n�	>�Z���������~�MUs �N�Er��xXc)O�%�~7Zz����&���#���ۭH���8�~���p�9�}��%Z3'�_��z�ӑ?jv���A�f�� ;$ؙ��v��������e���{�{���5(�����tC"-w�|���@���>��v=u�������6ghm�!=�y����h�}�BK9�H�.�c�T'9~�ʲ�GO�2o?�M��;]X��2�^WV���[%�c��\n$̱Z�)���2����_�*��!?9+�9D�s���J�z�3�I�犼C95^T�,+Ⱦ
� �AH���g���	�'�Wا[��������P3L!�F@�4%���V����*�qu|$z)��~�t}�Ft���i����'�,0��.b$ �([����
-�k�8���҆�|n��*�Y��p*Urq��;n��ra}�To?�M��;]/d^Bg�t��P	�x�[U���zy��<�hV�q��KPi8�����m��d�7������N\Q
7��0���Z�I��y�BR�J��?1;m�!=�y����h�}�#�?�G7�K��fC��t7V��eG�u���;��l)P�u��F"lܵ^��UŚ�p-�q��F@�u��w)�S����w����0~J�FI�n�w:Z�ZH��7u�Hߵg6{�I"H���cs}S�q��c7F���"wN��i��ӯ�0��\�4�s.)s:^�emߍu�M9Z�U����k|v� U�7C��H����b[/�<"����iN��{ ���Oz�-Y#дS����RRɤ>��y�m�!=�y����h�}����u*�V�xy�V��ݚc�rE�]7t۸�~�MUs fq�Ȉ��3RyE�'{_~�������C��.�Ė����D��&�$��(�X���I�ZV��W��x$���G��\�4�s|��Z�w��K�?g�W���7�:;�tp�{�k�7C��Hno��І�|�#}�{��N�Er��xXc)O�%�x��#y�D�+�N&	r�O��C��0���۞�^�n��t�r�}����r~%�w�>��S�C��ߊk'�4+.���`uI�[l٧cJ�^j�u��w)�S�3k:�(�-7��Mv�9\��(
�m�ó(��8�:r&@����p�T�c&�׸P)o�KӜ�u��w)�S�5� �p9�AE�t�ݙ����?g�歺4\�8O �L#Edɲ�<a6�}�%b�VJ #����ԁ�����`e�TS��\�4�s���rH
>TT	q��$6�0��2Y��-zX��Ƈ~�MUs �W_��i�~�����e�~9@�����k�8���҆�|n����{y��T���̦�=G�Tv��J�Й�m��C��ߊk'�4+.���`uI�[l٧cJ�^j�u��w)�SU��T�d�7��Mv�9��Nb'R��E�Kܑ�8�:r&@L���Qep��p�R��$���wT��xݣL����RL�a)=�y�~ ���H7���#h��@]7����7C��H��e!3֎�,��	�;�J�|(��jrHS�w�MH��j���r���+W��YJt�,�y"r� J&g~���c*& z�s�ђ�B�~f��0(�/��$ }2����T���Q���!i��ӯ�02�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vce��%;��I2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcN���HR8�p��}K��f<�,=K�F~�?|�[_X��ˆk�=�r���x�i��p�7��Xi9�
�ѹaB��Q�//?�s�m/C�N{a�9O!JoE'U�Y�y��
r�)�Y¹w����i��T!ix�AH�k[�^��_�)��6�$`Y���%�5�1�:�Ω�`<4}��)�Y¹w�yB-j&?��ј2��<��e�IC�_�\H�F?t�(����5�����~�Y��3g�ݜ��q�©�����Lu�m��+�����3�Χ��nEA��"0�qv+Y�y��
r�(����5�����x%~Y�1�:�Ω�S�T�;Ϗk[�^��_�)��6�$`���Uh7u+��T��٤�2[51g~Ӝ��ajƎ�c��(r���U�ј2��<��e�IC�_�\�����@J
A��w|�<��y�~/r�I��
����&�ɬ� VU+I���ť1k�`��'p�@�I�?g�f��m���6d��h�Ɵ�Y��FqqDt���,��B	hI�ˋ���Z�ZaPpJsd��E�#�ڊ<?@��[	J��;��2�F�P&l������ nU�IÙ=�H��[[��Vct�:��RE��Ok��@zL͊�q���Vǃ�����������-N���\�vņ�Q�]�ޝ��(��U��֜��3�b9���с�'sIP���1>y���Mw���1�Z���=���u*K6HT�����N��2�F�P*�7`����\Z��K���b9����4�6�t�8֩]=$����n�j�Q�ȧ��M*�'n�^0o��~+�ݗ����5�hbvk~�#x��܃Ae��'n�^0o`�U+�PAs ����
D�ZLN�	���b9���P9b��8֩]=$�?�R��n�~x�9̺��\�v�T?�7G|`^�R@Κ�2e�J�Pn\��J��H9��\�v�T?�7G|`^�R@Κ�2���C4�;��+���c�'n�^0o��~+�ݗ{,�
w��|ݔ�3�(n�'��b9���:&�>��sw�n���7[q�m�J�5�d�,W�� nU�IÙ=�H��'�PD�j�j2�%�5]��I踵}�=Ll�����&}0�@�͹ ��I�Q4p�/�;ϔW���1��ݥ�U� ���_�g)�X��Q�u������(�ʉ�I�,B�E?�xu����ma��u��ۯi\�q���Ìݣؤ	��#<��0a ӫ/��m�A0`��A��L�>�c'�'n�^0o���?��%%��XK���Π��yGb���u*K6H �i7�sp>ι��QG�����U��7�ܥ��2�\Z�ؿH�jGjh�rO-�<i���A���U��7�ܥ��2�\Z�ؿH�jGjh�rO-�=|-�e1|E�A�2����ma��7I�����5CS�|iɋ3���5�x�}+��U�p�[�����ma������	�I	"k�+���m l�o���ma��'f cTw��� +@���a
��|���\G�Y����-�,��Lt�2�tN�By3��<�]�!����M[��Ǣk/�z�xEQ�����5	���]���>����C���"����Y%T��BPe.��xu	�>��l%i�-\1��pz��S⏸[��c��Et�Y�{'%s�h�v���5���T�`�|��K�z�L;Л��Z�n��[��{_8�Y��=�}�Vݨ��������P���Qi�]2�y�Z鎬�����,�q�����CsYl���#�]�!����M[��Ǣr�x�e�X�����5	���]���c�A�L'��!�a��5�%]���a(􆿳����^��;�j����Y%T��BPe.��xu	�L$�����//��kOT$���]׽������E��@IE�U����S8����;(���5�%]���a(􆿳����^���#}�{�,�k,^+a�@IE�U����S8��$FW �9�װ?�p���5�%]���a(􆿳�ؖ��d�I�� �:&��I�?g�f��m���6d��h�Ɵ�Y����>3��w-iu�`���`�+N��?���&���#�{�0;�}����\Ҥ�Yk"1/��n5R�%�9��o�Dc�c~Ou�$�&�V��L��O��݄�$��F�Ճ����n�~8���a~�d��"J�A��S+e ���p�I��'�{��Ń��Dt�G_$�n�>߻��]H#
ZM��2 �єV��߼
�dgn�*�Q3#*�ۍc(yoy��Ŏh$���K5�!�>��y�P}��O��ꅽ52����$�Qu�&�<��G�JHn��z���z�O҈d�G}%��9��(��&��P��(*� ���Y�8 )�\�~xy��S��c��څH�8��)%sEW�o���開���?�`�7Ue�B �z��?�<W�$��Xo��Q��F����p�X��#�ڊ<?@��[	J��;�P4ǲ �x���\�E&��u��±�sR�{F3�_� ��0���c�B\����iW5�˦���X��lM��A( ����_�h3��{I��Z��H1�$ԠI�*U2��53��7�r޸��zL͊�q��$�%����#*�ۍc(y��p�r���C=2崝���v�+ʢG&q^�`
�c��><�$���|�r�HzL͊�q��C.W26K�~BvGޣkQ�A���ۖ��S�<Ԣ�E,�J�|R�ZLN�	��~m*�S%���^̽1��H����8�n�����ea�P4ǲ g�{�]4�W/S��8(�E���Kt㲎�������1#��Z�����XP��Ȭ���7���{r��bߣ$5/H�r�is�T�,�G��x�&[�ͧ�?Y;�L���9�D_�3���U_�+X�܄�֝���b�Bϱ�����7���{r��'6���;8=�g��U-�e���b P�G��x�&+8@V����L��\�E�V�6IWJE�r���秹�3I^�v�%j����L�de��-@��F~*7���&�_���/���l���F�8���/����RY��k�:A�	S�r��AR1<�N�؆�B��W+`�x�o���{��&�e�5
��Ib����rs�i�jf� l�Ǜ������CyW�f�tR�wX�����/��&����H���	N^�U��J��"ї�!~;��i�̥%�CvK���9u$d9�cx�S�����S8����ٺ?�R�^Ƒ����"X��[��Q[R�7�dט�w���V���Ĉ��r�]@Ԫ��d��ozL͊�q�����-���$�mo�6L���RY��D�of�7���A3�(N��㎏qló��|����=%+]Bo�A;h�F��O�i���Z鎬�������(���`$�P.eE���	fd�L;Л����׫�!�dט�w���f�ܗ��DX<�c>1K �:;k�+��b9������|L�K�)x�?{���x.�Knq	6�q�i�d�<om��'@�(��P�����k!� �J��/�oxW�}�zX<�c>1K �:;k�+��P4ǲ ��V �-�{q�������ތ�1��\�v�M��r�&�(vW4��`��?B��ž�'�t_� �e����Eck[�x�X��u�?�=�r�@^7&ģM�'n�^0o�<:�W�_�l�J;�RQ�y�� Y{q����'6���;8=�g��U-�e5/�=��kp�m~|��8yL2�����ތ�1��\�vŶ�T���Ĉ��r�]@s��I�λT�v��1���2���I��'�f�Nd+l��_]���T��\�vś��Z1`�x�y�Zglё�H�a)�r7�r��#[� B^�.�ߘ�)�I0M�/�s���'n�^0oPpkiq�o�H�MPq6.���fa���ӵ#yӛp�Tr�j.`#2��%0�$��Xo�U)+N���l~�U��tb@�s��\�v��/��v\�?� Zh�R������A^�7
7��Pt�e'J��\|YX�<I@1���t$I+�V�6IWJE�r���秹�3I^�v�[�9q�Y�{'%s��.|Z�����8��''6���;8=�g��U-�e5/�=��kp�m~|����U0��{ �=�%����|�r�HzL͊�q��C.W26K�~��^̽1��2������j{�-`VpN'O��h���]���!E����z���Jx�հ7$�K�2g�(#�.+ ���"��|���it	�TU����z~+Yi=��o�IÙ=�HVkLs��dJ�+���LQ�{p�uR�R�W�u���_�)�Y�5����`KIR*�fN����ތ�1��\�v��|z���m��P���ݪ��*h���'�aM�l��S�J*�Rs�08�b(�� ��˽��r�Q�gL#A=��a��'�-�O�Y�I�4];ˍH�P�(e�X�+��it�D(�	�}�]�O�hf>Ŋ�)4ԑ������~��7����g�E�����&��Z�4��軬P��|AC�JV�f}.�Б��+�B\zm�x�R���-�a3�i�a�>���t��.�Չ_:s�83���;�T ������]�W\(���;AD�S�/xm����r�in��oK=��\I@�ZJM)����d�8��⺞=I߀%)�	�b|s(��dט�w��]a��1qh_�n�To�[�C��-��JHn��z�Lqܳ<��J*�Rs�08�b(��E,�J�|R�ZLN�	��iԹ�08�@����gGNc�&�Ia�΁�a�n��!�`�(i3�n`5�fK�\w��0]b!��u��ܼ��	�!�`�(i3!�`�(i3�d�٣��c�A�L'�}g6��gf�Nd+l�Yҽ֗��i�ܰAb!��u�9*�"FP>����!�`�(i3��c�SD釛-���>T��`�z��Y��),�B۸��L� s�j8����DzL��k]m��6(�eZ�W���D��g�[�$��X�՚��l��Hr�<Uee�N�����H�OM��`�@����gGW�RJ����@{2귑��?4��44�|�%�|>`�|��K�z{�x���I�
�ݴR����,D�+�8��io�iA'R�	:�@�F����?�S��I��a\Y���};l�-��;a�������q�f@����DzL�����A@#֫��/�*ܑe�W����n�4�`t��D����M����A�m�(%�$�p��9C���1{Ģ� �z��^-j8�b!��u�ϟ��7�4Xe ��g[���
��D&e�2l��4(�de�QV踫g(�r�N�ǁ�f�TpD��ZOUi3�|)sՀ]�N��&��L�t��n�����!/��A3�(N��㎏qló]�b)�L�uf�Nd+l�Yҽ֗�2�0]�J}�
�?�a���k�_د@�CP�hWpH7���
I@1�ؠ&���Z02��`�z���n�j�Q�,���B�L� s�j8 ��*���v��W5�+k&v�IzZ鎬����
C��8q��f�kN�ı/���^�"�k'	-��>5i�[r�~s����R9Y�}��`y����@����gGKCYb,�q�K�M3�gwe�ŉm�m�jp=�>��o�
�v�ξ���I��RhF���t�>�˞1�����NR�^Ƒ����"X��[��Q[R�75�e`��9��əS\��O�=�Q���d�٣���������ݹ�0���f�Nd+l�Yҽ֗�)�|����P�%.^F�	��lC��U�T�\ ��Z��| �Ɛ�
�CӞD��m�q�/����g��d�٣��c�A�L'��!�a�~s����R9Y�}��`y����@����gG,#�g���b��Bg�� ��x��ό���.�}�
�?��:�,��mj�(���>����׌7<���������	N^�U{xN��i>r�<Uee���R�}vJ^�k��76����,Dk|q��K>�X$��V��ƇBHx\�'���Xw s4S�'�i��`�z����k!�\Z��K��uk�)�~s����R9Y�}��`y���h}Nw���Tc�~y��i�v1a{J�����u_7s�9���on�-�6��
�jW��D���M���o�G�m�?E]Gƃ	��[�x�X���+���LQ���"X��[��Q[R�7ݓ��E�/�����H7��[`���"�y���[�ͧ�?Y�f�kN�ı��U��+�Xa�H(�˕-+��B�Gݓ��E���vj��$ƇBHx\�'���Xw s4S�'�i��`�z����k!�\Z��K��y|��!k�R�^Ƒ����"X��[��Q[R�7ݓ��E�?\(8�e�!�`�(i3	r�&B"K�͢'����&���Z02��`�z����k!�\Z��K��^�7��u"�@����gG�Be|�����p&"&��MN���OON�
_�n�@/%{�;����f�kN�ı���}J�|���|���=�|�������n9��g�剤_��<��d�٣���������ݹ�0�������Dɵ�p�AJ�e�$��Z��7T�ߘ�)�Iƃ
ᾆ�x�T�\ ��Z��| �Ɛ��B�D�F �(����C�EPj�x�Z鎬�������(������t�\~ �g8Yw���k��$a(􆿳�ټ*w2�56��B�D�F a�^��D���Q]� _�rs�i��d�	�6%�����ׄ����ӯIJ ��`y����@����gGD=�^�(+�o\�FO�Z鎬������_�,���t��h~>#���d�٣��v_���Zo�ݓ��E�ȸgG�
��U,�(�)8���0y�	ű�;<9a�A��Y&��v�8:hJ�tV�nQ�rV{1m�V-���"X��[��Q[R�7ݓ��E��~>H���U,�(�)8���0y�	���T�<�2h�^Y�=R�wX��}�
�?��YN
��)e�3ݓ�V�?�f���,(���B���̴_��EI?�R��n��am�Za(􆿳���2����.�ɷ������5ʦ�q��T�ٮ|�,
������|�FIsŭf�ҿG�p�PR��{�&�8���/����,D ��Hl�E�ɍ�rH�ZAԢ�a\��F�dH��|c_�m��ġ��,�z���a�R�wX��}�
�?�����|���3ݓ�V�?�f���,(���B����_T���a�aq���E���ss�T�\ ������q�f@[�=�5x�.��Ӄ�7s�9���o��S8�/ #O�)R�^Ƒ����"X��[��Q[R�7����n9�jsrCm�k��Q]� _�rs�i��d�	�6%�����ׄ�hNݽ!�q�
�Bk�i�����B��' ��`y����@����gGC���yK�E����FZ鎬������_�,��T:���V�b߰6rh<xZ��j�
����d�R�wX��}�
�?��Pۢ����зq8�Ј'���Xw���,DH�v����ܹ����� �]�!����w�Հ�x9���7�.�I�A��7s�9���o>��l%i�-�u��Y'G-+;X����Jn,���`ό���.�}�
�?�ʬw�S��]+W��L��'���Xw���,D
zds)�
��g��#hi#����0z�cUL�J=��'EّD ����R�^Ƒ����"X��[�d�a�4$�b!��u�G9�:Q����v�z`�!�`�(i3q��T�ٮ|�,
���]�x}NI0���ԏ�.fOe	��q��"o��Q[R�7�)�`E5�j�W����+G���tJ]J�a:�xZ��j�
�iB{�Z�_�1�����\�H��/Sg�w��'o�D�P�E6���2����.JL���Z'#y�>�)L�����#3� n���a�x���w�K��r�]�4�P�l��=5;�<��|��k�8���/����,D��ǉã1X�v1a{J�j�f�At�-�=ѐn[���0y�	��sC宸I))����A�m�(/!���La|#9���b!��u�p��j����l�,9��!�`�(i3q��T���E@~����`y����@����gG�`����1�#��d_!�`�(i3ғ�vq�\[$Q��
�̞��>�_9�R�5;�/�O��� ӫ/��m�QP�*Hd���"X��[��Q[R�7�����bp�WdM4@��z(��e���b�ȵ�ixUS��F�dH�/�O��� ӫ/��mo��7�^�1�T�\ ��i3�|)sՀ*�şxˏ1��o\�B/��'����^\����b�Bϱ���w�K��r�]�4�P�l��=5;�<��|��k�8���/����,D����y�[�l��姹�g�YӅ:�y��Fp����L�de��-@��F~*7���&�_ƃ
ᾆ�x�T�\ ��i3�|)sՀ*�şxˏ1�iA'R�	��}E-�Z.��0�W\[$Q��
�̞��>��b��v݋N��������(($��R�wX��}�
�?�K�\7}�W,��+G���gÎק��-y|�$i�PiB{�Z�_�1�����\�H��/Sg�w��'o�D�P�E6���2����.�>��왩��k]m���E��Y�W�������a�x���w�K��r�]�4�P�l��=5;�<��|��k�8���/��%G��lyp1��>��kQ���� �^/s�1��p�E����F�f���,(���B����Ӝ$��BS�>�!/�_�n�To�[
MQ9�F�D�P�E6�q�l�.iAb!��u�L�Y}śT�!�`�(i3!�`�(i3O�=�ͦ����Jg�Z�n��[�]�u��yb!��u�[��m�U�H"҆>X�b���0��q��T��J�s���
�k��!a�tc�&ck��°������R�wX�ո@����gG��l��`�°�v�z`넥^�?�úAV�!s���0y�	��sC宸I))����A�m�(};l�-���~�]ݟ�R�wX��}�
�?�K�\7}�W,��+G���*�1S�@:8��=�?I®|�,
���]�x}NI0���ԏ�.fOe	m���h����$�'	�|#9���b!��u�[��m�U/|w~S."��|	�WI�U,�(�)8g��dT�W/S��8(�E���Kt㲎�������°������R�wX��}�
�?�K�\7}�W,��+G��ܼ��)�@�ғ�vq���q�41&q^�`
�c��><�$�X~��\��o����׋��`y���h}Nw��������j𛚆z�Ji��U,�(�)8���0y�	�z��SR:g()��ikp���H���F`���G���`y����@����gG�:,Z�g�YӅ:�q��T����<�սѡ��`y����@����gG�:,Z���@K�]�q��T���~��]�{�NլU]��g��U-�e,%�0g����Ed��>�^�v1a{J��8�P��Ά���0y�	��sC宸I))����A�m�(/!���La|#9���b!��u�}c��ko#a��|%GP"G�wk��r)��ׁ�a\Y����+���LQ���"X��[�d�a�4$�b!��u�G9�:Q��F��P�?��ě��+P"G�wk�١��	;qS�>�!/�_�n�To�[r��}k:�~�ȧq�6a(􆿳���2����.JL���Z'#y�>�)L�^b٫
z�����㞣ɐa�x���w�K��r�]�4�P�l��=5;R�ˊ	183��r`AZE�T�\ ��i3�|)sՀCeFJ5x�_�k]m��5L5@�m��R}>&_B�\[$Q��
�̞��>��b��v݋N������M}Ĭ���1����X�[��`y����@����gGQ��6��'�֤���n���6����?�& �.�|�,
���]�x}NI0���ԏ�.fOe	m���h����$�'	�|#9���b!��u�G9�:Q��Y���6#HA����P"G�wk�١��	;qS�>�!/�_�n�To�[r��}k:�~�ȧq�6a(􆿳���2����.JL���Z'#y�>�)L�b�@_	�][�����a�x���w�K��r�]�4�P�l��=5;R�ˊ	183��r`AZE�T�\ ��i3�|)sՀ�6�S2v}�k�����U�n޶���^.�]�|�,
���]�x}NI0���ԏ�.fOe	m���h����$�'	�|#9���b!��u�}c��ko#�gX�o��"�,�>E��P"G�wk��r)��ׁ�a\Y����)���8˩��F�{a(􆿳���2����.0��jOT��.m��K�+���w�7��'�b���b�Bϱ���w�K��r�]�4�P�l��=5;R�ˊ	18)Dg�|4��`y����@����gG,#�g��C�x!�H�g�F��'�ey�u��iB{�Z�_�1�����\�H��/Sg޶��j�}a�cf�g��U-�e,%�0g��սÕB\�6N �S���}me":l�ny��Fp����L�de��-@��F~*7���&�_���/���l���F�8���/�I����"�Oi9L�:�k]m����.aQ��-��b�Bϱ��R<�����á�~O��L;Л��|#9���b!��u��Ɔ ����;ƹ��:iq��T�ٛGS�����n���㬺ƃ
ᾆ�x�T�\ ������q�f@�]�gv���J�����_�U*��ө%�Sg()��ikp���H���O�=�ͦ�١��	;qS�>�!/�_�n�To�[
MQ9�F��g��U-�e,%�0g����]�gv���J����k̇���APߺ0��A���ۖn�a8�O�=�ͦ�١��	;qS�>�!/�_�n�To�[
MQ9�F��g��U-�ez�r�6JL���Z'���V��H?Ә�%"Q䛚�z�Ji�!�`�(i3!�`�(i3!�`�(i3зq8�Ј\[$Q��
�̞��>��b��v݋N��������(($��R�wX��}�
�?��x�������E��0�Z�7W�:��G�z㤧{��B��+ H!�`�(i3!�`�(i3ȵ�ixUS��F�dH�/�O��� ӫ/��mo��7�^�1�T�\ ��i3�|)sՀCeFJ5x�_�E��Y��Q�
w�8D�t�%o�V�g�yl��6T�T�D��ao.\C�k����-�|�,
���]�x}NI0���ԏ�.fOe	��q��"o��Q[R�7�)�`E5�d�G`5[��{#ŸFn�H�~M�!�`�(i3!�`�(i3!�`�(i3�E����F�f���,(���B����: ��ao.\C�kHgN�����`y����@����gG�7�{�mo5i,�Ĕi��)���!D�����ӸI))����A�m�(!�`�(i3O�=�ͦ�١��	;qS�>�!/�_�n�To�[
MQ9�F��g��U-�e,%�0g����]�gv��JeYSWe^E˔ �y=k�2�u���F�O����!�`�(i3!�`�(i3úAV�!s���0y�	��sC宸I))����A�m�(/!���La|#9���b!��u��V3���L�瞩w�j���@ΙN�[���-ل9�#c�ᜂl��=5;i�
;G(ɐa�x���w�K��r�]�4�P�l��=5;�<��|��k�8���/�I����"�CeFJ5x�_c(H޵D�ҏ@n�ɒ�[��iB{�Z�_�1�����\�H��/Sg�w��'o�D�P�E6���2����.JL���Z'#y�>�)L�����/s=s��4�+��_��A5W��v�8:�W�]�IVt���0y�	��sC宸I))����A�m�(};l�-���~�]ݟ�R�wX��}�
�?��I�_Pg<���7�*w�ɝF�l�u�*Ha���J*�Rs�0��7n�����a�x���w�K��r�]�4�P�l��=5;R�ˊ	183��r`AZE�T�\ ��i3�|)sՀCeFJ5x�_�k]m����DބiM��ө%�Sg()��ikp���H���k�XLF�iB{�Z�_�1�����\�H��/Sg޶��j�}a�cfC?�Q䨈��Q[R�7�)�`E5�j�W���yͧT���E��UH���4�������=�?I®|�,
���]�x}NI0���ԏ�.fOe	m���h����$�'	�|#9���b!��u���j�4��k]m���k�����A5W��v�8:���h�|!\[$Q��
�̞��>��b��v݋N������M}Ĭ����s�������Øf}�
�?��I�_Pg<ˉJLg�2'�r�G� Y��vrk�;}�f���,(���B����: ��ao.\C�k�ף�D�~�z$��8���/�M��%�p@!�`�(i3!�`�(i3>�3x̪�1�]�gv���{V�-_8���G�7W�:��G�z㤧{��FJ��iB{�Z�_�1�����\�H��/Sg޶��j�}a�cfC?�Q䨈��!&��F�!�`�(i3�mJ�0�6�b!��u�G9�:Q����D����1�Q�
w�8D�t�%o�V�g�yl��6�������	��oT���0y�	��sC宸I))����A�m�(};l�-���~�]ݟ�R�wX��}�
�?�����4R�ت����¿'��x!5����z�Ji�ȵ�ixUS��F�dH�/�O��� ӫ/��m�A0`��A���q_{}�g��U-�e���B�/!�`�(i3�mJ�0�6�b!��u�I	�����g[�s6{޴�i��)���!D������eW�d/=�y�H���|�,
���]�x}NI0���ԏ�.fOe	m���h����$�'	�*��/qRrm�ڨ�hծ�)�`E5�R(R�X���Ǹ���m�(��k8һ��6����^.�]�|�,
���]�x}NI0���ԏ�.fOe	m���h����$�'	�*��/qRr!�`�(i3�p}8�JL���Z'�����5qo��o�����&Sq�aj(��;���Q�y�QF����V��e��a�x���w�K��r�]�4�P�l��=5;R�ˊ	183��r`AZE�T�\ �ͧP?��;��$��Xo��4�!`��] �v"����W=D��'n�^0o2d���or_�B&��p�)Y����2����0/ܤ�(g��V아�nu�����.>mP��=�]:�J*�Rs�08�b(��n�� ���'�̗����#!d�+I0���ԏ�.fOe	��Cja����.)۞O��\�H��/Sg�w��'o�;��ވ�H��=#+��^n�r���n�(D�G�\ϫ\ʃ�1�9M��p����=j����s̓O "*B�^�b\��{��7���	(k�t �j�&.U}��le5�`���pɷ)A���	��s~d�0�@�W�o���{� ����i9v1�#��d_�U,�(�)8���0y�	���w������(�xk.��:�9l��"X��[��Q[R�7�u��Y'G�D厺��+/s�1��py��Fp����f���,(���B���Q��ǺΕR��ӟ-��ҫn$��_�n�To�[�d��WB���Q�n��-��`y����@����gG�!��V�B���.V��:��^��[�@g�#�ڊ<?@V��_?i89��c�[��GR�D^;d9ךp�+�n�)�o��Ca2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�/�����D"��K��(q�8�(�7yv}�!�P���Ħq�e�����<zA�iKF5����@��~˼��N�ǁ�f�T�ka%���:w�`�w5�O�%E#P�NK�z�R'cf����e�u�Vf�Nd+l�Yҽ֗�	����s*;��|B���r������*!��?�d���&�LS1c�0�2��$c���EyE-&�K^�G�u��0����.�����w���,��h����h���D�ҏ�6=������|���x��@��ǀ�D=�A���ۖ��S�<Ԣ�G�nJ `G�p�P�i�����;��|B���r����P���x�NS��7���ڙ�Q�Ր?!�`�(i3����;q�V5VM�dj��;q�:5A��p9�{�Jj3ų�z���_ΩI4��欱���j���1#Y�p���+�ϸ�i�	��+@f�Nd+l�Yҽ֗��x���`�;b�-�2�V��	��y�U}'FS��@	�<����2��EVA�ڦ�c4V�o��&���	M��3
�v�v-}�	mpB(p`D҉�Y~�y����u{ᵿ������6�~�5�O�%E#P��1�<������D66��~p�=m@�<����I�?g�f&:��r-,|�C�}�M!�`�(i3t�iZ]XF�hx��G��!�`�(i3��x��&^�B�wj$g�X;p`�ct�:��RE3z%�u�܆!�`�(i3�����ݱ������]�`�g()��ikp���H����>�#P�'�̗������צS0��ݚ�Н����8��T�h���}둮j\����C��rR#K�p�ݚ�Н��K�^��Q��G�S>\.�!::tm�0�i.�9!�`�(i3eX+��f J�"e~��O��!�i�3���j�\�"����ݚ�Н��� л�|�9I����o�u�/!�I=�+��2Y��kک�x����y���ݫ�ф���F�)!�`�(i3���ȍry��	�B�'��a�F�,�U6�Q�L��!�`�(i3��0�&�ͭ�U젩`#�4>?� �1!�`�(i3��"����M몴PBoT�ݚ�Н�?V��j�c�
���!8ϟ��7�4�Mzuf�?ǉ�=�2��}���zgm##��V5VM�d6��0]�1�v�9��s->m�9V��Vv��8>�=������iG��Ӆ�+��T�����D3���Dc�c~O�ݚ�Н�R�7h�,b0V�u�Q�ݚ�Н�¥������]n��-��w¹��<d�,��L��!�`�(i3��.��֞�������i�-�;8|,��3
�v�v-}�	mp�S�\�/H����8��p!E�t�0f�?ǉ�=�D�&��� �4V�H�%p"��R0�]|$�f�?ǉ�=jo���po�h0�h�#"
s���
|�1�0j�!�`�(i3؟��)�`U
]�,J��)v#��������6f1�W�`t��9��V�9<�6�Q=3���~�ǝ�,^ajķ�ʡ.>�!�`�(i3�2*Q=F���q/���<�����7
!�`�(i3�dv��oTN֢&@��&!�`�(i3k/�z�xEQ���*[UxG!�`�(i3��|��p��PIQ#�C,0�?���!�`�(i3��9��稕�a�/!O�f�?ǉ�=�2��}��CϾH�)�V5VM�d|�v�W��I4��欱���j����H������!�`�(i3q�\E��0�]��8ƹ��+5�4��c �&A�5I��RhF�� ��*�C�Js��I�HN��R��?�d���&����J=R���v�Q��/����T�m��+���J q.GJ����~s���^����p� 
���n	l��Q;�im��ȍry��	SƏw0�������_ۧ�-@t�/�W/S��8(�E���Kt㲬��MK�L�zg��p��I7��-5l*���T�I7��-5��5Z����+�t2�0�趦����'���o���a5��2Y��kک����Q��K�葀������Q��K�1#V���<��+qѭ�+g[�!�`�(i3�R6BQ�A�J�e�!�c�A�L'D�g�=a�iA'R�	9��&�f�ݚ�Н��w,�������-����rs�i��5O
T������Q��B%��߿�	G[4���$�wӨj]h���կ��~Z�V5VM�d�x�8�� ��ݚ�Н�{k�h�+��4�%�|#�r��8����AO��!�`�(i3�ra5�k�K�s.�֡mh�l�Rk�X��a!�`�(i3��3vS�vN��%u���ժ*)xJe��hy��)]W��7#OOJd֯�y��j��k����U{8�C,0�?���!�`�(i3E�l�����5Ƈ���	R����
w���Q?1\B�@o��[ea�8��������?9|[�,HJ
?�?J��k����Lt�iZ]XF�hx��G��!�`�(i3 k��v(�Âv����Y���a\Y����+���LQ�f�?ǉ�=�]V�H7'�R�^Ƒ���)ύ^��R�^Ƒ��f�?ǉ�=j:�Mpp�}�(�-lc4�j
Թf�?ǉ�=��X�u��
)\Y����4MT2g�ȨQ�?�Q!�`�(i3���ȍry��	SƏw0��П�+�
8'���Xw�j�7��9*�"FP>���뭟Q��ǺΕ�A�m�(�]�	��B7Ԅ��SƏw0�����.>H'���Xw�j�7��9*�"FP�jV�$d,H�Q��ǺΕ�A�m�(�]�	��+#Cxz!B��2��}��̏A��?�ϟ��7�4Ï�6]S*�N�ǁ�f�TpD��ZOU	XT�1�wӨj]h�z��?�9��V5VM�dn�0�I4��欱���j����,X�|H*!�`�(i3u�l�T.��:��]]t�L�t��n=蛗�+N���������$��+#Cxz!B�`
 ֢����oC���b�J
�g��*�7`����\Z��K���䈷UJ!�`�(i30q���Q�L��!�`�(i3bs��2[������	�;�ݚ�Н��\�LtF�/�X�h��E�i�m}66j�"Hs��ˑ1Ms�����x����A@�Q��ǺΕ�A�m�(jj�*y��}�+�ϸ�i$x���z*�7`����\Z��K������]NS��.�g3Z�j5�{�ݢ��e��[њl����{O��c_`J��Y��)�.����ߤ��/��5�O�%E#PP���x�NS`|.^~�/W�/�#+*f�GR�D^�-�����6j�"Hs��埏���7�VL%�ǅ�����xF�~B�@o��[ea�8��������?9|[�,HJ
?�?J��k^"�u��.��������֢&@��& k��v(�Âv����Y���a\Y����)���8�w�A���k|p��z~�I7��-5l*���T�I7��-5��5Z��S��ك6
��^H��sp�]3t�ҧ{����Q��K�葀������Q��K֭�B������t��˳3[�u8��R6BQ�A�J�e�!�c�A�L'D�g�=a�iA'R�	:�@�F���m�6�&Zt%��m&<�jQ	)>_Z鎬�������(���ڔ6�.���Vd��\_�>�� �?"�Q?V��j�c��99�)b�+5�4��c �&A�5I��RhF��F4#_�h��霧�`�x&�e��A�:��]]t�L�t��n���%�(�N������	\k�`��B7Ԅ���ra5�k�K�s.�֡mh�l�Rk�X�Q��ǺΕ�A�m�(It8Z�QC�P�v	��Y4]:C�2Y(���˜V�Q��ǺΕ�A�m�(It8Z�QCf�?ǉ�=I��
�[��b=���|��p8=�[Ǵ��p���@Z�|�)՜�4�vIn�������23�,�M(���������b�8�dX�↨q�©�����<��p����Գ+ڍ�P��o�|��S�x�l��1:�N�*�x�w,�����<v���G�=���Q{�1�a-���7a
��r����~v��f�?ǉ�=ct�:��REvє�&���ct�:��RE3z%�u�܆j:�Mpp�}�(�-lc4�j
Թf�?ǉ�=C��[�����p��@LC��[���Ը��q�������ȍry��	Y��'�����0��"��S8�TkF����v1a{J��bC������
&0$o�<������N�u��]�!��	Ǹ�y85��U�z����@{2귑��?4��44���u1�E
�2��}��̏A��?�ϟ��7�4Ï�6]S*�N�ǁ�f�TIX����B7Ԅ��3�kM�}��s.�֡m�\�&e���Q��ǺΕ�A�m�(D}����4��2��}��M�p}��ϟ��7�4:i�P.j*�7`����\Z��K������}�4%6� �7�'%��e�툙A_�u�N�ǁ�f�TIX����B7Ԅ��0q���Q�L��֭�h��O�"Ԫ b]�4>?� �1�\�LtF�/�X�h�����]�]�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vczңh��p�^g����>Θ�Oh$d�I�v|����3��8�>�o����f[o��X���u%�RAo�������s�_c�Vr���J��:���闩R��M���'HY-��Yk"1/���]���lw]�찝���n	l��Q;�im��ȍry��	�����ň���)��a�<P��C�*�7`����\Z��K�����+��g�]V�H7'�R�^Ƒ���)ύ^��R�^Ƒ��f�?ǉ�=߼��� ������iW����<5�;���?$l7�z!�`�(i3R�c4!`��������F�)�_�������� "5�]�/��@��e:$h�7�cl.�	�C˟B�'��a���r�N��(�����������c�����:��IK��<��"��4�#:S�.?<a���k�_g������rVu,� �C?wm��:S�.?<a���k�_�aY��|rVu,� �{k�h�+:S�.?<a���k�_�~v� 1���\�9nW���z@]c�'���Q<��dq_҂T�q�w���I4��欱���j����%�`:�����Z���F%�X�ԃ]�����Ձ�=�n�4��Ǳ߁R�^Ƒ�өwo��Z��Ac<�p{�5�O�%E#P��"�=�X���?�`d�!g�lu/��g�)�I��#�r��8�3����Iӷ��}Dq�f��.��.f�Cz瀿3�z���]�D��V5VM�d��?s[�rY�C'Y#�6�A�m�(n$�(^i��$r�t�}iV��	��y�� �P�qN�h���w3&�D�U�2Y�û�gj��EYzȧԡ�/$a��F˯�+)Ƒॉ,����g��U-�e a⣃_B7�}�!��a���k�_]���^��m���PH�F��׿]=ͅ�J<v�z�����	�.�g3ZrZ�0m�\�n�8�Z�Ѽ)E��J�V�6j�"Hs�l��J�&�E�U�P�)��ꬪ1�7��/z*q+6j�"Hs-kS�Y�n����P����z4x��x�L�FZ�1�.SS�Zs�c<�^<�H�W+��W�*%b;���`,9�H�W��`�z��Y��),�B۸����H�V�7�}�!��a���k�_,&�BV��̷_��yC��S8��(�RJUlJ�,>�]y�P��l�}0��]T�o8b���L-kF˯�+)Ɠ�E��G�6��J{�a�Ĉ��r�]@�l��}$�SK�mBqJa��ߛ�����R�<1�V��	��ylK�;���aT��3G?�d���&����'-*�!�Fr忒@2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc���߱QD��G�����_�����o��A5D������1φ��<�6�@a� ��fFMqlg{y����i�q,?5q��r�I�	s�<�e��BFbs��2[�a��o���H�RtV�^��j�4��݄���K7͍��|��W&":����@|����^a�nu4Bޗ��jw�	���|#HK��=�O�-v�*_�mS8<�n�ݚ�Н�G��-�HG(l��l��n�]�!��	Ǹ�y85���]��^������.'ӟ�X#�r��8��vJ�F}��I��RhF��F4#_�h��WU�~�F˯�+)Ɠ�E��G��;b�-�2��;�P�t�5$f��_Ub���uQL+��φ��<�6�h��^�`��_���w���;2j�X�&_ܑ�Y(�����&� &��( a⣃_BR���Bk�d0��jOT���b�S]���o"83��Jn,���`�rs�i�Q�*NެC�T�\ �͜����Ƀ<;0V5���yʟ�SlX(�(�y�Vx1h��-:.02�v�Կk*����]�a�m��rÏ	��f6���H��\���
y���%~w4�( ����@����y�|M�rs�&
Q�j+�B��,"b����<pb/�yn��]������JD}����닓.�`�3��.S����l[�Te�H�qfP�0���@f��HG�e�#in4~������^����lWw6�b5�/
X�y�b�O�lnO���u��m���P����H�!��(zfx�q�Q7��f_����hѓ���Q�Y���\�'Zb>���C������];h�/�c�{��lq��:)�
�9LeQp�K�}q^J=��ڥ����Ⱦ
��7t��i97��EN�Q,�SGŹ닓.�`�3�^��D�Ϲ܌��!��!�`�(i3!�`�(i3!�`�(i3.[�Kδ9~��q6g�yF}���V6K�K*g�B�w���	�e���0��Qܓ'{w#/ B!�`�(i3!�`�(i3!�`�(i3}Y;�jns->m�9V��y��{�"���b��Bg<���P�5]'\gWg��	�Z�kfc?�#	*]]�iI9�o«IX0F�M�bw,���b�S])ެS��B�H����Qw�c4~Nr_�mS8<�n�ݚ�Н�G��-�HG($R�i�Yl-ۼ��%�ۙ�b�S]���o"83�C�
���W����Uh1�b_X�XV�b�z'hۉ)��d�7�qĹ߆�p�h��d��JXl'�T��~��Uг�|<!�`�(i3e<�Ia��la��o���H�RtV�^c�{��lq��:)�
�9LeQp�K֣����[$R�i�Yl-H�1O�N�
��2a� 硙�t�\��j�4�<�..�4��xu*���Y{�<���^�[�-l�H�=��
ڨg��U-�e�,���6+�HN��R��bP�63Z�t��Ě����E�i�m}6߸��S�Ȍ��7���9��j�4�<�..�4����9q��e��b�S]���З�}ߟ�r�Q��b��Bgk"������m�q�/���e���W�.�]ؔVG�A����}������݉}]%'6̳�ه4�tZOuLI݀����j�R��m�q�/�Wv�A��F!��D�����k$ !�`�(i3!�`�(i3�T�T�y��~yZ�|	����7i����S�y\��&�+������e����y
 <]9�(b���J��:����'X��u�>�
��`��<�
�d�ξ���Ix���Ka�0e��_�:��d���!i�wӨj]h�}�������IЫ�Is�8�w\�PPO�s"�6
���}Dq�f�����,�ǰ�|���]O_U�In��u�.�g3Z�Ǵݵ���{ �4"-��Dd>�STV��	��y�N �T�Jə�?Uhi+�h�#�����@���"�v6�z'kKǹ|���|u��R+��O�r!�J��:����G��-�HG($R�i�Yl-�x�f7﹏!�`�(i3�I����~u/��kOT�:�,��E�O˅!���U��+�Xa�H(�˕�3�,�Oj��j�4�q��_N��¼��=Bg����@N��ޠ����u�Y�KG�ξ���Ix���Ka�0e��_�:��d���!i1�����j�QXv�5���P!3)T짤.��.f�� D�_\HN��R��?�d���&�(���o{ٔ|0����T�4(���;��|Bh��� ���H���-��Αo��p2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc{�-���鏈wƠ�q����V-l���`�qf���?v�q�2�_:��p\I��� �W�G��!?�d���&�db�\EXP-7�vqq��I�?g�f��r�F�5��I^ξ��ݴg��S�ZCw]�찝���n	l��Q;�im��ȍry��	^�R@Κ�2���eip���,��x�y�ZglZ�(�SڬG�ݚ�Н�3A��gd�J�`���nU�gF�r�f�t���MK�L���NK�3�Fq)~�@�&-)���(`��ү/�O'�=��k�+9=�]V�H7'�R�^Ƒ�ӭ�i�\�>&�&i��&�C�/S��ك6
��^H��sc4�j
Թf�?ǉ�=�t���\�W+�[Z����4��#o�C��[���ԗ��6%�ac��� �G�T(e���ZYM	^:�x�����:��uL�e����kn4@Q�/�!�`�(i3�5?�&P-�C7z���Ɔ �����Vd��?�+�p!�wӨj]h�jsrCm�k��b![笐��vj��$�<��RN��B�'��a���r�N��(�����֭�h��O�"Ԫ b]�4>?� �1�������c�����3
]!p�a���c
��X���(� ^��D5�|أͽgF"?�Q��ǺΕo�G�m�?a"��-K8?�d���&��D�U�2Y��2܌�B�ja�M)ikZ!+�[�x�X���+���LQ�wo��Z��Ac<�p{�5�O�%E#P�G�dE�h�k]m��,�۞��	���B�è������iA'R�	op|��G�E�i�m}66j�"Hs�ĖYS�������P���w������x��	A�V��u�Vx�%Ls�N
�u�}�T�\ ��;��|B���r�����N��t���[���mt�\�lO��cb>�g�D�I��)���W�w��fD�g�9��,Y��(c$�,w�R���y���,!�뱁�c
��X��u��V�H�t����M~V��	��ym��θN�,�2#��2��{�Na{Gj��J�1	�<������UG���{b62�tstJ��:������L��t��*����	��#�����.�g3ZJ���V�)��w� �1@�`�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc:#�c>���D��ν������4����6S����'HY-��Yk"1/р�{:��'��F�N~Y�}n���t�iZ]XF�hx��G�����=�-�o&l������g����=�tt"���O�����J��a�U"�������o��\�l�Ϧ���I�:뼥<7.��H�ʱˡFZd6�o�·���~X�~���$^!!�`�(i3uwТ�
2������}�k�+9=����Kp&�@���k��-��w¹��<d���	fd,���9^-��כ��p܏�<
DN��X;p`�Vx�%L3z%�u�܆��O���R�^Ƒ��!�`�(i3*bL�(R��u��n�k|p��z~���8��'@���k�� tZ�u���ߘ�)�Ij;��q,��
4#!���ڃ�"�!�`�(i3�������t���ck��,�:�N�*�x��0�&�ͭ-��i�m�T�੝�hy��Q�#<4^�>N0Θ��;b�-�2�>c��?Ӈa�/!O�f�?ǉ�=�<��>��%@��4��).i���SRX$��V����覭L��G�dE�h�����?�O̀���vj��$��覭L�q�\E��0	ozqPx�6_s/��g������n3�x�h�k�t]�<Lz�l#�V��H��<�C�Ar��� f�Nd+l��p��;z�_��s�֙R���Bk�d*e��\@8GS��`n������ct�:��RE�QS����>�wo��Z��Ac<�p{�5�O�%E#P�P����9��g�ܧ*y*J�X�$����aV}�������,���1����,H/������,�ǰ�������'����2�,bxqX��g�9��,Y�����9C�������u8q��ǵc��5�%]����8�B���ow_;O
�J��:���闺����ő��"�\�!�{~����DKY�����|f���+X�E�k?�i2�.[W�w��fD�g�9��,Y��(c$�,w�R���y���,!��HC�d��g���'N3 �zY]�埅�t�į��>�n��-�U4��\w��˪?�-�l~�U�n��(���_��s�֙R���Bk�dNmyM<�G�ۺ�Ub�!�V��u��i�_:�����k��$�8�B���ow_;O
�J��:�����A��AC�m]���z2�nFW�JyS��f
t斃����u_�*5o]E�HN��R��?�d���&�c�����|�� 7�G�Yw�R���y���,!��HC�d��g�[��f��*�)|/P2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc:#�c>���yn�4^4 ��#�$G�l����M���R'),��`ތ@�'��|0;��|B�v��䣞�a���~�(����5���&<˴m���q~�i���}n����ϸ��#|S������3[�u8�~6���q���)�� �tNU�:|��6/��������рӚx�f�?ǉ�=����Kp&�@���k�֖sK3��!�Y�7#�xI���E���v:ι�Y+W���F�^�Y�7#�xIvє�&������0/�e��9�SW�Ty��5!�`�(i3���0/ܤ�(g��V	QY��K*�+W���F�^��NP&�2�������ȍry��	��0�&�ͭ-��i�m�T��!�`�(i3k/�z�xEQTl�������l6��\�LtF�-��{����"�2��}�������Ə:S�.?<ߌ�LM�a$,�۞��	�rVu,� �{k�h�+-�����*��$�q�ʋ�b�Y�S�:ԫL�S��S���ONY 
~�F�,���XF:6/��������рӚx��^�̷ؠ�ۈ`4�`�����w��oe��7�uvWދ�qc:_U)�<�&#�+���LQ�wo��Z��Ac<�p{���`�2�G�Y���s+��6�.'=��!�����tAC��g��op|��GKW℀4ٜ���,�ǰ����������^k�3���RӒ};��|B���0�2u��[�탓��t����M~V��	��y<C�.���@6��[��C���D3�N*��ј�Q��O�بeD�I�,����y���Z��FkH���޴�ik]���7�i�s+��6�.m���1�Μ���,�ǰTm�v��G��y2Z��Zk��Αo��p2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc{�-���o���sp%T�a�U��M�u@x���m��+e�(���n�JŬ+�|�C�}�M�ϸ��#|S������3[�u8�ct�:��RE��]n��xj����R���it	�TU����z~���MK�L^�R@Κ�2'�̗�����b��Pp��h�5,Wlr�r%)cA�&�C�/�h��=;�_�8V��F�x)3پ������ׄ���MK�L�P�i2s�4<��!I��5��4]�폮h;e��w�5�ϟv�BA�IH���O,8(�6k�4d�Lt�2�t�U젩`#�4>?� �1Y��
�iC�&8�,��Q�L�������!�`�(i33��(b�W���5�.SƏw0�����98[Ɯ��X)�:O̐�V2XUt�{#	�x�=�tneX /*;63��dn��AmOeTky�q�\E��0</���/�u�[-�c]^�ʎӦ�V�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}�Y�o��}�����k��h`�H�MPq6.�yܤ�܎~�J���^W�������������_�ft�m-���L%�o5j
�^q�&Ѣ�� ��&6�%�@��n{�\�<:���\���D)�g�%v�=̽�0Բ�ȁ��;�<�h�kIp�#J,i�~X�Z�o�x��o��ײ]�4�Kq%��M�Vr���J��:����;�	��o�g��}>�IM8e�׸J�q��G��m��+�Ƽ(��h�Dc�c~OPM�^-q�x�l��1:�N�*�x��
[N<p�U��֜��3�X;p`�Q�%�+2�j;��q,�?�Ho2��ݪ��t����$�fC` ��\�H�MPq6.����gQ'�|ݔ�3�(n�'�f�?ǉ�=$(��>��������	���i$;��|��T�.�l�.θ��q����k��,�:�N�*�x3Lv	̅���X;p`�(�����֭�h��O5�tx\s�l.�	�C�
�:qEp��:��Z)�"r��^&���贵[�л���7#���=
 �4���ߩ��ݚ�Н�p�n���d�)bU��� �Y.�.�g3Z�7�4��~��=�>�:|]η��E�<���5[�������0j|�~{b62�tstJ��:����s͟;)f���d�jO)īIX0F�MV�ҁGG`5:�����8-|�D�H����Qw�c4~Nr_�mS8<�n�ݚ�Н�+��%�k<a�E�Rq���my$�N��o�/���;�Ra])n#���^a�nu4Bޗ��jw�	���ݚ�Н��}�АR�38v�s3~�0�����&G!�`�(i3+��%�k<����m��5vȹ|b�7�ݚ�Н����F��O��;b�-�2��;�P�t�5W?�;��@qz�_vrrL�����^�%�P�m�V��	��y�f�HYs��uF��82�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��OC�0����t��[���P��EC�`�/�t�KV*�3?�|��T�5�d�,W�He�!� U����z~/�}��j,NJ��:����8���SY�N�o��C�0�_E,�8�o��_�Rv�䩲$��GQЌJ
�յ[+8����"sS<�0�zG�������&G�wӨj]h�(%����K7͍��|��W&":�;b�-�2�k+Q�h'�Ȝx�5W ��̫(� h�ҩ�-��)'�E��ȷ��#o�]�ʄǾH/�d��_�mS8<�n�ݚ�Н���4�*BqC��~�;ϔW򻐗�NGq���ÌZ>u�,R�� h�ҩ��wӨj]h�(%����+�uB;y���O�	���lC��U�T�\ ���:5A��pfĉ>99��A0ok�ª���l��������t�|ݔ�3�5�}�]�����nv��~���$r@H�RtV�^;�jmT�#��|�!�[�w/	��^#��4,�Q��+�uB;y6R��*Q�z�ׯ�1p1�Z���=��,�����!���2�(+�uB;y���O�	������v�h��4y��ij��X� 2!�`�(i3>_�Bnˌw/	��^#��4,�Q��+�uB;y6R��*Q�z�ׯ�1p1�Z���=�1�(�yj�!���2�(+�uB;y���O�	������v�h���ў�L��-����!�`�(i3q�\E��0����G�t���m�� �ݪ���CyW�f�tR�wX��!�`�(i3�	��x��ݚ�Н�����l��q�P�oV4ʐ�}	�[���&�ŁHL�U���W�����&G!�`�(i3�wӨj]h�(%����Z鎬�������(���/%Z�ڄ^1�B/���q%U����z~(����(]�U����z~)���	6�!�`�(i3�Ra])n#���r����!�`�(i3�� ߌ��̷_��yC��S8�>c��6/{v=~P0:Q+�3yK������v�h!M�T�ĥ��P�7� �:5A��p!�`�(i3���F��O��ݚ�Н�fĉ>99��A0ok��
�:qEp�;�P�t�5
�:qEp�;�P�t�5fĉ>99��A0ok�׹�3��܌o��oŵE=�[�P�X;�Z��;_��8W�w��fD[�P�X;�Z<0)��TG䟳��LQ�%�+2��k��kK�I�Q4p�/Cj���C�1A%^�Q��U����z~/�}��j,NJ��:����8���SY�N�d�}����U��)���Y;e�iK!���d.O.C��|#HK��A(�c���_G��Hb� h�ҩ�{k�h�+E�g�������(ӈ���m�r����̢k���F�KD�Vr[/}>5��0�B� �b�Ъ���l���{$����^V���!ֿ*Y��b"���LQ�/81tSjv��wӨj]h�(%����Z鎬�������(���[���-���W�6?��jsrCm�k#��2�bD�=�^݊��}Dq�f���Ě�����}Dq�f��5ߧE4��HN��R���IX0F�M����m#p��ܸ2߆X�.�g3Z��S~����l�I�k2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc:#�c>�ϓ'�al��p;��|BB�Q�ˇWv�A��=a��0� �Jeh|�*�7`����\Z��K��7�,�B/�Q{z�
wb����T�}ɻ*�7`����\Z��K�����6�~�5�O�%E#Pe�6&	 �|��k�|��SSB������a�v'�m����o��_�Rv�䩲$��GQЌJ
��`���φ��<�6�15���Dl=*�QN������"sS<�0�zG�������&G�0�9&،�j�W����+G��ܒ���7�_
�uz!:�X	��sC宸I))����A�m�(mq?��qU�՝� s�#0�ʂ�j�Ï��	�l�lM�3 H�RtV�^܌;���d��-��!C�� R�Q�&�2���)x�?{���x.�Knq��5+*��d�@���G�X���.��ġ��,��5+*��4br���qP�V>t'�̗�����F��~1tSjv��0�9&،�j�W����+G����v�9'�͘6��q���j�W����+G���|��nZ����ݚ�Н����F��O��;b�-�2��;�P�t�5W?�;�끣�os�鮊(=�"v��Iw�6!e�C�7ª6��J�����_�U*��ө%�Sg()��ikp���H����c���鿉�X+�kQ��v1a{J�i�\��ou#�m ޶&�hbvk~�#x��#�H�޼QE1��v1a{J�&���e�� տ�:
hbvk~�#xo�������Qטg�u2]c
j���l��姹��*�ɿ�4J*�Rs�08�b(���,bxqX�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�ᾣ4��LG9�:Q��Ĵ��ޯi�-Qq��Pn9a�Fc��Ǔ��K��v1a{J��blv�Bo��"~6���aq������n}L�I))����A�m�(�l���q�b��v݋N�������H��YTN��r8!�k]m��
ae���K���c����P7E����k]m��GTH�<�g()��ikp���H����7�����\�H��/Sg�w��'o����̜�I0���ԏ�.fOe	j�)6)-
2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�ƹ9��PdG9�:Q��Ĵ��ޯi�-Qq��Pn�����G�v1a{J���!<�*Ha���J*�Rs�0��O�@�n�M?��h�k]m���E��Y��m���+)x�?{����}9��|�G9�:Q��Ĵ��ޯiڼ�ze��>տ�:
hbvk~�#x�<\��-��4�1���~!�`�(i3!�`�(i3!�`�(i3N��r8!�k]m���E��Y��m���+)x�?{��
0#`�1�������f�l��=5;�B�uʡ ޼QE1��v1a{J����%]+a�����G�v1a{J�&���e�� տ�:
hbvk~�#x+[.Sk�NA�I�_Pg<�l��姹�n4'����3
�v�v-}�	mpJOv�����o\�B/u�:o+���	�����aq��c�:X��Wwl53�e�'{w#/ B!�`�(i3!�`�(i3!�`�(i3G9�:Q����v�z`���ө%�Sg()��ikp���H���R����� ӫ/��mt����� ���M��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>h�wbk�$�޹���M�,!hޖ�A$�P������5d�������y�:Fa�7���W"�P�K�0_f��3%�:��IY]��r$ɓǃl[�Ƶ�1tSjv� #��zG���J����(�u���p��,\���͔5��:m�\�H��/Sg�w��'o��Lͷw���]�x}NI0���ԏ�.fOe	�ߣ
����Ra])n#���^a�nu4Bޗ��jw�	���ݚ�Н�y�}�6f&r#o�]�ʄ�g�s���������J*�Rs�08�b(��h�P�\�䖬n���S滑����ZLN�	��;�uO��Bu����aGl��Z����pG�p�P�$�c76u��r��M�yx�,�G#y�>�)L�Y�S�:3�g(���27:։�X+�kQ��v1a{J�c�Q$ a�3��}Dq�f���Ě�����}Dq�f��5ߧE4��HN��R���IX0F�M��uR�Y�A��-�R�͢��n-(�p��Kث��@�uj���V��H?Ә�%"Q䛚�z�Ji�!�`�(i3!�`�(i3!�`�(i3�I����~u͘6��q���j�W���]�B� �Q�ސ�՝.�&J�m�(��k8���0[�d�G`5[��{#Ÿ�&Sq�a"��ř�!�`�(i3!�`�(i3����;q�a�x�G9�:Q��Ĵ��ޯi�^�0��ͅ�a��;���=����qFq�w�鎷�Z,����d�G`5[��{#Ÿ�&Sq�a���y*/@(�_��%$>_�n�To�[�pI�
K�x�������E��0�Z�7W�:��G�z㤧{�̌�͚�3�_�n�To�[���9�P�4�D�pc�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�2���$H�WdM4@��z(�ﳔ$@PJ+5*�轓�A1�J�����)����Ҿm�(��k8���̜�I0���ԏ�.fOe	���X�a1p��j����Q�9�|`��Y�m�k?j!�`�(i3!�`�(i3!�`�(i3�a�x�]c
j���%��g:������	����^,�:��O�?�I))����A�m�(!|�α+���s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc9g�O��B~K�\7}�W, D�cg�}ŷ(K���}�;]MBg2Zr�G� Y�ҹnЭ:��#�@����ۭXX���E��O�;]MBg2Zr�G� Y!s!��xlJeYSWe^E˔ �y=kt��w��X����xQ�1���~!�`�(i3m��i�*�JeYSWe^E˔ �y=kAu5��ݞ<\�H��/Sg�w��'oD+���4Yʁ���Mյ��#�@����ۭXX���E��O�;]MBg2Zr�G� Y!s!��xlJeYSWe^E˔ �y=kt��w��X<���H1���~!�`�(i3m��i�*��9$��i�Yi䚠疛!wFii�v1[���b��v݋N�������(X��#�@����ۭXX�WŚl��E�d�G`5[��{#Ÿ�&Sq�a�"Ĝ���$��a�vw����~m�(��k8w��?L�@^?���W��j�[O����k$ !�`�(i3��䨘J�\mo5i,�Ĕi��)��ۺ��fyd�F�O����!�`�(i3!�`�(i3(*�O�q�@��i)&
�k�����oT`kz��9$��i�Yi䚠疛!wFii�1�В���,؁C�*&#�4?�o�5�h�B�ˊ��6Ԩ{�1{&��� )S���z�d�G`5[��{#Ÿ�&Sq�a���y*/@(�_��%$>_�n�To�[B���v��؁C�*&#�4?�o�5�h�B�$5z&�D�� ި�6v ӫ/��m����	�����tj/�Ս��6Bj�!�`�(i3M�yx�,�G؁C�*&#�4?�o�5�h�B�$5z&�D�� ި�6v ӫ/��m���l]�f��EJ,�G7```+�ֶ������x�������E��0�Z�7W�:��G�z㤧{�r�(��mo5i,�Ĕi��)��ۺ��fyd�8]|Fl���1F#�֞q�F����&U;��]�x�'��x!5�kz���[hin5�҇�?�b��v݋N�����-
#?�QAmo5i,�Ĕi��)��ۺ��fyd�e�՝*U�޸I))����A�m�(^?����8������k$ !�`�(i3�~�7p����nt=:�+�_0c ���a�vw����~m�(��k8!�`�(i3!�`�(i3!�`�(i3׾ŞWsuz��"]c�#y�>�)L��H"҆>X�(JdT�ݙڈ�KK?B�&�_j�	�Ȗ@@��x�������E��0�Z�7W�:���p*�h<��I0���ԏc�r�(����I����~u��a�vw����~m�(��k8un��7� ӫ/��mt�����N��r8!c(H޵D7W�:����p�A�B��+ H!�`�(i3!�`�(i39a�Fc���M똡����o\�B/�u���a�x����r͖�k���$,�C�7ª6�JeYSWe^E˔ �y=k�2�u���e�՝*U�޸I))����A�m�(9�*��� c(H޵D7W�:����p�Ǎ�͚�3�_�n�To�[���9�P�4�D�pc�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�2���$H�WdM4@��_�U*Cw�Hm���9��N	{8G9�:Q��Ĵ��ޯi�3>٫F�?��"��II��jÇ+�_�n�To�[
MQ9�F�GM��QО��i/R�c� }!�`Uc�gC�!�`�(i3!�`�(i3!�`�(i3�a�x�]c
j���l��姹� �p�B���#;%%�.�4����
��\�H��/Sg�w��'o�֕ߝԀ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��4?ڇ���WdM4@��_�U*Cw�Hm����a�vw����~m�(��k8�����9�Xy+�Mk��L

�F����&U;��]�x�'��x!5�kz���[h�b��v݋N�����-
#?�QAmo5i,�Ĕi��)���!D�����ӸI))����A�m�(^?���W��j�[O����k$ !�`�(i3��䨘J�\mo5i,�Ĕi��)���!D�����ӸI))����A�m�(!�`�(i3�����wP?��i/R�ce����� .����mo5i,�Ĕi��)���!D�����ӸI))����A�m�(�[?;$�\��E��0�Z�7W�:���p*�h<��I0���ԏ�?��Ds�-�w���+kGA��ݼ��r����!�`�(i3�o�5��!<��y�@�v�&Sq�a��z#׊;w�����f�l��=5;F5E�]q�hf��EJ,�G7```+�ֶ�����rS����u�}�Q���GM�о٫�o�}Z�\Q;]MBg2Zr�G� Y� {l��	�:�f�?���tj/�Ս��6Bj�!�`�(i3M�yx�,�G���V��H?Ә�%"Q�ܦfM� �L�Y}śT�!�`�(i3!�`�(i3G�&ց�*�p8�Iט��ō�Zm\�l��ì�A���V��H?Ә�%"Q�ܦfM� �'9�5���c(H޵D7W�:����p�A�ԍ'8����J�������"��<��y�@�v�&Sq�aj(��;����_��%$>_�n�To�[B���v�쟎��V��H?Ә�%"Q�ܦfM� �in5�҇�?�b��v݋N�����U-�pë��";Yy\'{w#/ B!�`�(i3޼QE1������m�(��k8һ��6ݕ��wp>�\�H��/Sg�Al�a�;�����9�Xy+�Mk��趵��1�F���������m�(��k8һ��6�D��)��	u�}�Q���GM�о٫��s�~�L�1{&��� )S���z;]MBg2Zr�G� Y� {l��	�g�yl��6T�T�D��ao.\C�kT���/T$ǩ����m�(��k8һ��6ݕ��wp>�\�H��/Sg�u-Y2�G�1{&��� �5掼�s��ݚ�Н�!�`�(i3K7͍��|��W&":!�Fr忒@2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�l~�1��n��+��o�JJ�tsq��T�G�'�q��;��y�-���2���澝ߚ���PC� �ˆ��*2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�WOtl��[��m�U����#3T��_�[g���pj������e�S�[�k]m��
ae���K��ʭ�!c����fx'v�ao.\C�k C�Mh�n �O`�Ag��ۭXX0���?V�#=uz��ɜڈ�KK?Ba���$_��v�z`��E�4ki��w�K��r�]�4�P�l��=5;���o�1g��U-�e'+]�{0C!�`�(i3!�`�(i3!�`�(i3AԢ�a\�g.��m6]c
j���%��g:���1nSpɃb6vJ�pZ� 4�F�Α��Bʏ,�:��O�?�I))����A�m�(�UVh�hP[�t��#��l��姹�xAQ�Y;x����$����7��=�S:t�L)��k]m��l��e b6vJ�pZ� 4�F�Α_)'!��r���U�4�8�v1a{J�j�f�AtT��_�[g�����,��WdM4@��_�U*��{��������
��\�H��/Sg�w��'o�GM��QО��i/R�c� }!�`��8
|�Kvb6vJ�pZ� 4�F�Α�v1a{J�j�f�At╔����̞��>��b��v݋N���������L+-�8���/����̜�I0���ԏ�.fOe	pۙE�����WdM4@��_�U*��Wc��V9a�Fc���M똡���iA'R�	s��]C�m�(��k8�4k_ł�k]m���E��Y� ,���� ��̆���M똡����o\�B/�u���a�x����r͖�1r����X�N�SF�vb6vJ�pZ�t���%�Q���� �^]�y܃fs�A���5��Q���� �^/s�1��p����;q�Zܑ��B$�䪜Q3N������2(wUF�|��: ��ao.\C�ktg����U��pqo�}9�-�_����NǨQ�~�^��>}�;�D#��2~��vNOgۈPM�r�]�4�P�l��=5;,��'ٕΖ�%����%2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�w�u��[�wbk�$�Z��Ջ`,9�H�W��`�z��Y��)h��{��Ķ�,�����F�!��cܦ���ҧ�v1a{J�)�3�� E!�`�(i3!�`�(i3�I����~u[��m�U�tV2�8�.�`��ai���Q��B%W����˩I4��欱���j���1#Y�p�� �VBD�!�Ĵ��ޯi��:��:̹��.�g3Z�7�4��~�U��{��0��L�r:h]��Ve.*�QN������s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�WOtl�ܨ$�`V1���cЉ�M�$@PJ+5*�轓�A1�J�����)����Ҿ���M���X���̜�I0���ԏ�.fOe	j�)6)-
2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�ƹ9��Pd�V3����C��z���Bf���a�x�G9�:Q����v�z`���pqo�}�;-�]�̓@?5�M%jWhC䨛��D)��C�V���3������G��������M���X�����9�;]MBg2Z�ܱ�Q3�!s!��xlJeYSWe^E1��b���t��w��X����xQ�1���~!�`�(i3!�`�(i3޼QE1���������M���XR����� ӫ/��mt����� ���M��2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�cRq>ha3@��[/�������ܦR'cf���³5��*�7`����\Z��K�����5�O�%E#P����ҧ�v1a{J�"M�X�m�Z!�`�(i3!�`�(i3�I����~u}c��ko#���uT�.��=�F�@{2귑����|�kI��RhF�� ��*�C߇���t�k]m���E�i�m}66j�"Hs�@��C�,ԭ}3Y�Z��E��3?�d���&�Û=�������fo��ZpW4%"������k�I��RhF�䂔�R�D����M���XH {��u��]'\gWg��	�Z�kfc�_	�Ƽ��S�J\7!c�2����X�G[��7�癆cgQw�c4~Nr_�mS8<�n/�"����5=��)Q���nF���<�W�.�P�	��
�Q�}����g�Z��3��a���!@�f")u��r��܌;���'����u��r��#�աl����aGl�97��EN�y�JB���PY~�y����o)�T*�c�Q��Ne<��t��y���'j��ݚ�Н�i#\��u�vc�jj&��G�9m6�̟�1��"~6���aq��3=]��m�D��-����!�`�(i3px!��ia��T)�
���l�K�>�������Ra])n#���r����`
 ֢���̟�1dN�<@Iv��nt=:��:5A��pfĉ>99��A0ok��fĉ>99��A0ok��$f��_Ub��7��G_���;�P�t�5�׹�ն'�U;|�� �R�SBJ���z`�3ޕ ���t�T��?E-h��`f���sd�G}%����3f闶P���`�3ޕ �7�癆cgQw�c4~Nr_�mS8<�n/�"����ZRR���dN�<@Iv��nt=:�$r�t�}ik+Q�h'�Ȝx�5W ��̫(� h�ҩ�y�}�6f&rG��Hb� h�ҩ�0�p9zr��XƤ5_���"~6���aq��k�7� r��H�?�k ���50f
V��.ᬵy��f�'XĘ��L�F.	-�L��&PY~�y����o)�T*�c���-/a8!�`�(i3닓.�`�3E�g�������(ӈ���m�r����Ra])n#���r�����+��9,(ZRR���&���Ɗ3I5=��)Q�]� ���_�hbvk~�#x��	���"��]ap�~��q6g�yF}���V6l;�<��'�̗����Ep� �����4br���^��D�Ϛ�-����!�`�(i3�N(	I��^� �&����	cS�6�=P�ݚ�Н�$f��_Ub�F�S�1 �$f��_Ub�F�S�1 ����F��O�}�	76�&�� Ӗ�t$�)�vxִ/pJ��#��p,m��Q���M�"/���h|����6�o8:4�I���c�90��G��6�iI9�o«IX0F�M��uR3��%<�X�7�癆cgQw�c4~Nr_�mS8<�nQ'݀�=�Xy+�Mk���[��9�my$�N��o�/���;�̢k���F�KD�Vr[/}>5��0�B� �b���H�����Yu�������&G����l�鞏̩jv�^������J*�Rs�08�b(��h�P�\�䖬n���S滑����ZLN�	��JFХ�B�9�4br���qP�V>t'�̗����S]�_�_��u��r��M�yx�,�G��i/R�c�'DV���b�z'hۉ)��d�7�q�՝� s�#���k$ �H�����4br���qP�V>t'�̗�����F��~1tSjv�!�`�(i3Q�>�H�((��"Jk�\p��j�������\�z�ݚ�Н�$f��_Ub�F�S�1 �$f��_Ub�F�S�1 ����F��O�}�	76�&�� Ӗ�t$�)�vxlP�6=��Nh�����x@�*�j��m�(��k8H {��u��]'\gWg��	�Z�kfc�_	�Ƽ��S�J\75�e��4��X�G[��7�癆cgQw�c4~Nr_�mS8<�n(�6k�4dFn�H�~M�h��,���ANʂ��t�Ǌ���z
A��Φ�gz(AٸI))����A�m�(��2M�`�̢k���F�KD�Vr[/}>5��0�B� �b���H�����Yu�������&G����l�鞏̩jv�^������J*�Rs�08�b(��h�P�\�䖬n���S滑����ZLN�	��JFХ�B�9�4br���qP�V>t'�̗����S]�_�_��u��r��</Sn���̟�197��EN��~�{�B��R��� �hvT�+]�x}NI0���ԏ�.fOe	��;csj/�՝� s�#���k$ �H����p��j�����8"c��"��]ap��e��>��Օ��qvdЧ^{�jMdGN���!�`�(i3��T��xW����˦G�m�(��k8��0�m���!�`�(i3�5ߧE4��!�`�(i3�5ߧE4�퉅�%>�rGO�D mWN��Ě���aT��3G�IX0F�Mm�(��k8��xh�j�W���5L5@�m�$R�nS�]'\gWg��	�Z�kfc�_	�Ƽ��S�J\7!c�2���j"�²O�i.����bs��2[�a��o���H�RtV�^G9�:Q����Z$�x$�֯� W97��EN�Q,�SGŹ�R���/�O��� ӫ/��m�A0`��A�2�����$r�t�}ik+Q�h'�Ȝx�5W ��̫(� h�ҩ�y�}�6f&r#o�]�ʄ�g�s���������J*�Rs�08�b(��h�P�\�䖬n���S滑����ZLN�	��;�uO��Bu����aGl��Z����pG�p�P�m������� h�ҩ�޼QE1��v1a{J����nFy� �����&��"]c�#y�>�)L�����/s=s�^�?��:5A��p���F��O�}�	76�&�� Ӗ�t$�)�vxģ��_�ڑ��� en��`��n5��=�8�`Lv�RU��n;3ѫIX0F�MV�ҁGG%4vkz����`���φ��<�6�15���Dl=*�QN����r$ɓǃl[�Ƶ�1tSjv�޼QE1��v1a{J���Ꭓ�[��^E4+у��b�Bϱ��b��v݋N������M}Ĭ��ʡ.,�-��̞��>��b��v݋N������M}Ĭ�����Gf�߆�p�h��d��JXl'�T��~��Uг�|<;�jmT�#�,l����?0G.{T�2��^/e��d]� ���_�hbvk~�#x��	���Ze2O�W.����M��p�#���F�H۷`"��]ap��e��>��Օ��qvdЧ^{�jMdGN���!�`�(i3G9�:Q��Y����(��U� P"G�wk��M똡��A�{�>�� ��
^�Mi~_�THN��R��bP�63Z�t�5ߧE4��Fr��j����bm&����T���Ꭓ�[�"�2�~�m�ek�}/�*��^��φ��<�6�@a� ��fFMqlg{y����i�q,?5qi��(.�j2��w�V�"xjzӝ���I(͂��-����N��r8!�k]m����DބiM�^E4+у��b�Bϱ��b��v݋N������M}Ĭ���՞)Ǭ�Q̞��>��b��v݋N������M}Ĭ�����Gf�߆�p�h��d��JXl'�T��~��Uг�|<;�jmT�#�,l����?0G.{T�2��^/e��d]� ���_�hbvk~�#x��	���Ze2O�W.����M��p�#���F�H۷`"��]ap��e��>��Օ��qvdЧ^{�jMdGN���!�`�(i3G9�:Q��F��P�?�u�$�+AԢ�a\�]c
j���(y�.
جH�)��
���z#��#��Ě����E�i�m}6O�D mWN��ܐ�}��s����$c���Dx<�Θy9����s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}�޼QE1��v1a{J����nFy� �_Y��t��3
�v�v-}�	mp����/�כ�"]c�#y�>�)L�����/s=s�1�3���3
�v�v-}�	mp@?��jV�H�I�_Pg<���7�*w�ɝF�l�u�*Ha���J*�Rs�0�ǳ7��y.+�F�$-�S:t�L)��k]m����\�6�=�r��J*�Rs�08�b(��g]�6��;b#y�>�)L�^b٫
zܫ5u�q��	�����aq��p�Rdae�Qטg�u2]c
j���(y�.
جH�h��p\��"~6���aq����{M�jX Kp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc������N��r8!�k]m��5L5@�m��i�*O����Qטg�u2�Tt$Ó6N�֤���n���6����?R����� ӫ/��m�A0`��A��7A�Ǩ�3
�v�v-}�	mpBR9ƭ�����fx'v�ao.\C�k�ף�D�~.8s�Z��N��r8!�k]m����\�6�EM?�ۄ�a�x�]c
j�����7�*w���Ǌ����fx'v�ao.\C�k�ף�D�~��pr����)x�?{���x.�Knq��!cI͸I))����A�m�(};l�-����׭�i�#�}��il��Rm�㭼�S}�S��S�C���+�%�t�*#y�>�)L�^b٫
z�.h��E��B\�H��/Sg޶��g�R6Ӹ�m ޶&�hbvk~�#x}���y���>��� ӫ/��m�A0`��A�;��ܞt�td���52�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�ƹ9��PdG9�:Q����Z$�xQ�RY�##�� �~�^#y�>�)L�����/s=s��4�+��_��A5W��v�8:D�!�̞{��L]Eц~_�֤���n���6����?��ө%�Sg()��ikp���H���]c
j���4���TS3���/k���m���+)x�?{���<m�N=-�w���+ާ�����ݚ�Н�!�`�(i3!�`�(i3!�`�(i3G9�:Q����Z$�x�vG��*Ha���J*�Rs�0K=X���d���fx'v�ao.\C�k�ף�D�~�Y�I���I�_Pg<���7�*w��D��q��� �~�^#y�>�)L�b�@_	���UH���4տ�:
hbvk~�#x+[.Sk�NA�I�_Pg<���7�*w�ɝF�l�u�*Ha���J*�Rs�0��|�_�Y�j�W����΂o�����4�+��_��A5W��v�8:'w/�'��γ~<����jVѭ@!�`�(i3!�`�(i3!�`�(i3 #��zG���J����0;�����5u�q��	�����aq��ɪw�*=>@\�H��/Sg޶��d��5��f�C�7ª6��J�������ߧj@QEM?�ۄ��I�_Pg<�(y�.
جH��O��U
hPߺ0��A���ۖC�#dG訠�O`�Ag�v1a{J�Bz��s�V��m���+)x�?{����}9��|�G9�:Q��F��P�?��4�+��_��A5W��v�8:'w/�'��γ~<����jVѭ@!�`�(i3!�`�(i3!�`�(i3 #��zG���J�������ߧj@Q�_Y��t��3
�v�v-}�	mpl�!����_�n�To�[r��}k:�2Y�ا 2'l:}��Q2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc]�&P��	��I�_Pg<ˉJLg�2'�r�G� YF��6�!�`�(i3!�`�(i3!�`�(i3����;q�a�x�G9�:Q��Y����G[�����a�x����r͖�k���$,�C�7ª6�{V�-_8���G�7W�:��G�z㤧{��B��+ H!�`�(i3!�`�(i39a�Fc���M똡���֤���n���6����?���$����;-�]�pR�$5iL�Pf8e���N��r8!)�5���sO���%�$�m�(��k8w��?L�@�b��QM!i�9�s��J�a$�Y �������G����1�E�AvY�5�h�B�c\��L̎C��fx'v�ao.\C�k�ף�D�~�Y�I�����s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�WOtl��[�t��#��l��姹�C�`N���$@PJ+5zqiS�Q#y�>�)L�b�@_	��}Pz1Z�ݗ�"��I�����f�l��=5;R�ˊ	18kQ����&|���BY��l��=5;R�ˊ	18EYx��*��O`�Ag��ۭXX�|ʡi�����Fz�!�`�(i3!�`�(i3����&���0���y�هj�W�����ד*(�os}�&à�m�(��k8�*�0�mI0���ԏ�.fOe	m���h�����̜�I0���ԏ�.fOe	m���h��֕ߝԀ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��4?ڇ���WdM4@�k̇���AEM?�ۄ��I�_Pg<ˉJLg�2'�r�G� Y�ҹnЭ:��#�@����ۭXX���E��O��j�W���bԽ�b��˔ �y=kg�������8�`Lv�RU���7xw���	�e��1{&��� �5掼�s��ݚ�Н�!�`�(i3]c
j��ʉJLg�2'�r�G� Y�)�?���I))����A�m�(};l�-��	}�<�Q"!�`�(i3�����9�Xy+�Mk��L

�F����8�`Lv�RU���7x�.9�?	��j�W���bԽ�b��˔ �y=kt��w��X<���H1���~!�`�(i3m��i�*��{V�-_8���G�7W�:��G�z㤧{����+c_�n�To�[r��}k:�>�hyȷ����wP?��i/R�c��;=~.�"�f!Hb�G����1�E�AvY�5�h�B�]�{���j�W���<�'��V�I�'��x!5�kz���[h�x�1W0�u]9�#�I���jVѭ@!�`�(i3 #��zG���{V�-_8���G�7W�:��G�z㤧{��B��+ H�ݓ�W���"r�DyA�S⏸[��t��7�M~G9�:Q����D����1�Q�
w�8D�t�%o�V\�Z�0��{V�-_8���G�7W�:��G�z㤧{��ԍ'8����J�����"�f!Hb�G����1�E�AvY�5�h�B�$5z&�D���ME�R�, �5��U���j�W���<�'��V�I�'��x!5�kz���[hin5�҇�?����XzR���bn�u]9�#�I���jVѭ@!�`�(i3 #��zG���{V�-_8���G�7W�:��G�z㤧{�E2p��F4F�[��\	.���#�"r�DyA�S⏸[��t��7�M~G9�:Q����D����1�Q�
w�8D�t�%o�V\�Z�0��{V�-_8���G�7W�:��G�z㤧{��ԍ'8����J�����"�f!Hb�G����1�E�AvY�5�h�B�$5z&�D���ME�R�, �5��U���j�W���<�'��V�I�'��x!5�kz���[hin5�҇�?����XzR���bn�������mo��jVѭ@!�`�(i3��dN���ub�z'hۉ)S���o޼QE1���Ꭓ�[��Yi䚠�5���u�L�!�`�(i3!�`�(i3!�`�(i3��c���鿉�X+�kQ��v1a{J���Ꭓ�[����$����;-�]�pR�$5iL�z#��#I	�����g[�s6{޴�i��)���!D������eW�d/=me�%b\%�I����~uI	�����g[�s6{޴�i��)�������T�\�H��/Sg޶��d��5��f�C�7ª6�)��%��+b�O~1��GM�о٫�S��wE\�!�`�(i3!�`�(i3�I����~u͘6��q���j�W���yͧT���E����ua�����\�ec[�U�b(l�rD��ЀUg]�6��;b�����5qo��o�����&Sq�aj(��;���Q�y�QF��fK�Ěk.�����GBz��s�V�r�G� Y� {l��	�m��ze��I))����A�m�(};l�-��o���n[�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcE���Q�K�\7}�W,��+G���*�1S�@:8S�C����0���y�هj�W����΂o���R��o�3��rD��ЀUR����� ӫ/��m�A0`��A�"��(ޅ���>��� ӫ/��m�A0`��A�,���$�n�M?��hS⏸[��א �k/ׇӭ��!�`�(i3!�`�(i3!�`�(i3����}>R� [�'a,�v1a{J��¸�k�Lpަ	<�%�;�ÇI���fx'v�ao.\C�k�ף�D�~���~�C9w��fx'v�ao.\C�k�ף�D�~h1��'�t�Kp(����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc����1 ��⒍~��Ĵ��ޯi��ŁO�(K���}�H[W2q�[�Kx�ʁQ7W�:���iޚuq6p��j����Q�9�|`ЉɁmwl��\�6��#P��Ѐ�5�h�B��ME�R�, m��
~�B�H[W2q�[�Kx�ʁQ7W�:���|���~�Fȯ+3�YE\����oW���";Yy\'{w#/ B!�`�(i3޼QE1���Ꭓ�[��Yi䚠疛!wFii��{s��ֹ�Em��r�~ʁ���Mյ��#�@����ۭXX���E��O�H[W2q�[�Kx�ʁQ7W�:���|���~�Fȯ+3�YE\L�}��鋿 ��
�Q�
w�8D�t�%o�V����������F>�w�γ~<�����6Bj�!�`�(i39<��`f�R(R�X���Ǹ���m�(��k8һ��6�R����� ӫ/��m�A0`��A�,���$�f��EJ,�G7```+�ֶ������]G��܎~:Q��z�˔ �y=k�2�u��܉�ӌ$/k�Bz��s�V�r�G� Y� {l��	�:�f�?���tj/�Ս��6Bj�!�`�(i3M�yx�,�G�����5qo��o�����&Sq�a��z#׊;w!�`�(i3!�`�(i3G�&ց�*�p8�Iט��ō�Zm\�l��ì�A�����5qo��o�����&Sq�ae:rmv�H�!�jT7|�`\%��u7W�:����p�A�ԍ'8����J����T"O5�`�7B��[�<?Ә�%"Q�ܦfM� �in5�҇�?����XzRL��MWX��DބiML�瞩w�j���@ΙN�[���-ل�{s��ֹ��!n)\HL�U���W�H�2^�/3!�`�(i3�0�9&،�R(R�X���Ǹ���m�(��k8һ��6��b��QM!Ϊu��U)�(*�O�q�@��i)&
�k�����oT`kz�)��%��+b�O~1��GM�о٫�o�}Z�\Q�R(R�X���Ǹ���m�(��k8һ��6�^?���I�^$D��Ҽ]G��܎~:Q��z�˔ �y=k�2�u���e�՝*U��eW�d/=4��b�Bz��s�V�r�G� Y� {l��	�g�yl��6����������F>�w�γ~<�����6Bj�!�`�(i3=��a���my$�N��o�/���;B����WN�Q���=�&�Φ�3h]��Ve.vrWB�i�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�WOtl�ܧG%�MP3ö�3���Cw�Hm���9��N	{8G9�:Q��F��P�?\��R?��f�I))����A�m�(};l�-��Y��bq7h9��n� I�&|���BY��l��=5;R�ˊ	18�׼�^`���s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}��I�_Pg<�(y�.
جH��O��U
h�07�;|''����˦G�͘6��q���j�W���yͧT���Ek�s���qa��;���=��i�uP=�z�}o*o���D)��ʱ�O�Ϸ(K���}Ǉj�W���yͧT���E��UH���4�����ˮ�N��G9�:Q��F��P�?��4�+��_碍�(H��(�K��k]m����DބiM�YG5`FFB���r����+C�ާ�����ݚ�Н�!�`�(i3!�`�(i3�I�_Pg<�(y�.
جH��O��U
h�07�;|''�)�?���I))����A�m�(};l�-��X;l_��Z2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vcq]�~��B�56e����bn3�qj]'\gWg��	�Z�kfc�_	�Ƽ��S�J\7������B�56e��Y�p���]nA(�c���_G��Hb� h�ҩ�G��-�HG(�b�'Be���0��_�,\��݇��h	��F���L��b��v݋N������M}Ĭ��ʰ"���(���B����: ��ao.\C�k�ף�D�~��(��ᩁ��@|����^a�nu4Bޗ��jw�	���|#HK��=�O�-v�*�Va�ir���M��2"���&�^��v�8:?�'��ᦾ�;���8���U�._�nQ�rV��q�t7�v�]��1���U�._�h�5,Wlr�r%)cA�r�(�%�pH�RtV�^��@�z]��C�x!�H�k��^)(���27:����i�k�G/�����	^%�R��^�Mi~_�THN��R��bP�63Z�t�5ߧE4��Fr��j������B�56e���D����a�.m��K�+���w�?�H$~��	�����aq����>s�P�T����ym) �S���}�cЉ�M1y���TJ*�Rs�08�b(����Ph���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vck�ss:mo3G��-�HG(�b�'Be�i�}���$@PJ+5y*���� �S���}�cЉ�M�V�O�SFl�A���ۖ��S�<Ԣ������f�l��=5;R�ˊ	18kQ����&|���BY��l��=5;R�ˊ	18�׼�^`���s�lI2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vcb��D�/�����	^%�R��aX��͟i8��m�q�/��v1a{J��U�Iv}տ�:
hbvk~�#x+[.Sk�NAG��-�HG(�b�'Be����\)Pߺ0��A���ۖ�w㌐g�߂.m��K�+���w�?�H$~��	�����aq��Ż%g�VƇ�m���Ar)���r����!�`�(i3!�`�(i3!�`�(i3��j�4��k]m���k�����A5W��v�8:C��4�I[��I))����A�m�(};l�-���j�	30�����Q��B%��>&ޝ�?1P��C&��b��Ɔ ����-˄�_-����dA�>�[E��1���~!�`�(i3!�`�(i3!�`�(i3-�E��%��v1a{J�a
�E��`���:�#�.��N�x%�M�RG�_`��z7{'#O�v1a{J�����ciA9*�"FP��� �mD��.1|��I�����V0�k]m��������fQ:b׻���3�v1a{J��bC�������N���� �VBD�!�Ĵ��ޯi�`͘�c�N&��H8|2�c�P�@��E�)�`L��%P��,���|�������[�i�*���1���"D���;�Ӏ�<qs��#�����M<E��'Z*)�?�R��n��h
:h����t�h��W+��W��v1a{J���&Y��V�Ԙ~q�9����t�T��?E-h��`f���sC>��Ӛ��S�J\7&���"�g72O!j���v�۲=�k2;�jmT�#bs��2[�a��o���H�RtV�^�G%�MP3�;ƹ��:i!�`�(i3��nF���<�W�.�P�	��
�Q�}9��?xs}�k�����|	�WIx����E2b�z'hۉ)��d�7�q�</Sn���k]m��D+_{6/ ���we��0�U+�qbp@�!�`�(i3[��m�U�H"҆>X� ��H�B�{_8�Y��=�}�Vݨ��}Dq�f��⒍~����v�z`��Ǖ��`���nF���<�W�.�P�	��
�Q�}���Mڷ��iA'R�	z�#,gB��3|v��Eb�z'hۉ)��d�7�q�Dw\����.m��TDZ��O$/ ���we��0�U+�qbp@�!�`�(i3�Ɔ ����;ƹ��:i����;q�{_8�Y��=�}�Vݨ��}Dq�f��N(	I��^��@K�]�!�`�(i3��nF���<�W�.�P�	��
�Q�}�k��^�1��dc�@c�����h��-����;�jmT�#�,l����M?��y�!�`�(i3�G%�MP3�;ƹ��:i!�`�(i3���G��x��?�S��K�+���w�M�7��<�1�����\�H��/Sg�w��'oª���#oM��:<��j!�`�(i3�G%�MP3ö�3���!�`�(i3���G��x��?�S��}�k���ޗb�Ͻq%(���B����: ��ao.\C�k�ף�D�~n��1w{��8���/��:5A��p١w��zj�v1a{J��湮��}6�/S� ����,��WdM4@��z(�ﳍ�f�_��S�>�!/�_�n�To�[
MQ9�F���"X��[�,�!���D!�`�(i3K�\7}�W,��+G��ܢN��_;��(���27:����7D!��%��g:���
A�%�q���F�dH�/�O��� ӫ/��m��M���	a(􆿳�3�m�
2]�!�`�(i3[��m�U/|w~S."����ʲ�P"G�wk�#�_wU|�1��v�z`넥^�?��F�dH�/�O��� ӫ/��m�A0`��Aw�zɝ8c��g��U-�e1�S������/��@���WdM4@��_�U*�u�$�+AԢ�a\�G�n봈2=��+G���*�1S�@:8M�7��<�1�����\�H��/Sg޶��j�}a�cf��"X��[�,�!���D!�`�(i3G��-�HG(�b�'Be��O����}ߟ�r�Q�C�x!�H��Yů�a��(���B����: ��ao.\C�k�ף�D�~n��1w{��8���/���}Dq�f��G�dE�h�k]m��!�`�(i3g��c���b�'Be���I-�X!�`�(i3닓.�`�3BڴQ��J�a$�Y �Mn__��q��ڍ$f��_Ub�F�S�1 ����F��O�}�	76�&�φ��<�6��'�al��p\ٿ�6�P)� &�]?�t�ϗ;��|B���?#�+Fz��Ԥ�Ԙ~q�9�C=2崝��tw�i�՗[�:X#x;2z��
�@h�5,Wlr�r%)cA��z>9�R��d���!i�6�5�p����M����-)O^��� �F��s]'\gWg��	�Z�kfc?�#	*]]�iI9�o«IX0F�M�v1a{J���&Y��V�scX{�X!,�'ž1�|�'����u��r��9��?xsTDZ��O$!�`�(i3x����E2b�z'hۉ)��d�7�q�`
 ֢���k]m���Ǖ��`�/ ���we��0�U+�qbp@�!�`�(i3[��m�U����L�F����;q�{_8�Y��=�}�Vݨ��}Dq�f��⒍~��Ĵ��ޯi�ʌ	���bS��nF���<�W�.�P�	��
�Q�}���Mڷ���o\�B/���2�>x����E2b�z'hۉ)��d�7�q�</Sn���k]m���E��Y�%��W#<e��0�U+�qbp@�!�`�(i3��j�4��k]m������;q�{_8�Y��=�}�Vݨ��}Dq�f�W����GTDZ��O$!�`�(i3��nF���<�W�.�P�	��
�Q�}����FYs96j��
!�`�(i3x����E2b�z'hۉ)��d�7�qĹ߆�p�h��d��JXl'�T��~��Uг�|<!�`�(i3e<�Ia��la��o���H�RtV�^9��?xsTDZ��O$!�`�(i3�i�<�~�y�j�q�7�AԢ�a\蟴���P`��ɠD(c!)��w�K��r�]�4�P�l��=5;���o�1g��U-�e1�S�������6���2[QvA�LO�>��
�I����~u�4br��
�uݟ�x��?�S��}�k���ޗb�Ͻq%(���B����: ��ao.\C�k�ף�D�~n��1w{��8���/��:5A��p١w��zj�v1a{J��湮�ձ������r���IbW�P"G�wk�#�_wU|�1��v�z`넀r?&��AK��sC宸I))����A�m�(�QNȮ���k/��m#��}Dq�f����Mڷ��iA'R�	�yvc�]k�i�<�~�y�j�q�7�AԢ�a\�G�n봈2=��+G��܇�c.}M�$(���B����: ��ao.\C�kf��_@Z��T�\ �͆�v�9��</Sn���k]m��������fQ�qr�~�룺���aGl�k/E΋*U���7D!��l��姹�C�`N��䍬f�_��S�>�!/�_�n�To�[r��}k:�d4��f��a(􆿳�3�m�
2]�!�`�(i3[��m�U�H"҆>X�\2�~|G��YN
��)e
�����z%t��#-�v1a{J���!<�b�Ͻq%(���B����: ��ao.\C�k�ף�D�~n��1w{��8���/��:5A��p;�x'_|~� �S���}me":l�n�������r���IbW�G��-�HG(�b�'Bep�w�{�̞��>��b��v݋N������M}Ĭ���F`���G���`y����ݚ�Н���nސ�Ѵ����-VL!�`�(i3��DKY���k]m������W�!�`�(i3I8�ѐv2zigzA=v)����;q닓.�`�3��}Dq�f���Ě�����}Dq�f��5ߧE4��HN��R���IX0F�M�v1a{J���&Y��V�kcZ�Z�f��;_��8W�w��fD��e���WƂ�\���O�!2ɵ��w�o��'�R<l�K�T�}�̖˄��O��r��'������ܦR'cf���³5��*�7`����\Z��K��qb	��G��W+��W���fy����φ��<�6�@a� ��fFMqlgd�G}%����3fEa�F��x��A�Z����r$ɓǃl[�Ƶ�1tSjv�-�E��%�k�Vx3G�)P<�ܓ�Y�Ra])n#���^a�nu4Bޗ��jw�	���ݚ�Н�y�}�6f&rG��Hb� h�ҩ�-�E��%�k�Vx3G��Mn__���ͥ
ݐ����%>�rGO�D mWNHN��R��bP�63Z�t��ܐ�}�Ea�F��x�j���NC�V��	��y���B��у#Y�wP-�H1�m��d�7�T
u�/%F���J���rG[Pt��H {��u��]'\gWg��	�Z�kfc�_	�Ƽ���8|bs��2[�a��o���H�RtV�^�Ɔ ���Ve��˅�E�g�������(ӈ���m�r����*qA����6\�4�@�� �-j�1tSjv��
�t��T&���LQ�/8"��]ap��e��>��Օ��qvdЧ^{�jMdGN���!�`�(i3�p�8H���v1a{J�ikl(rco��(`��ү/�O'�=�CyQ�/Ap�H�RtV�^�G�dE�h�k]m��Cw�Hm���Ɔ ���Ve��˅��ԝy'��Ra])n#���r�����G�dE�h�k]m��Cw�Hm��K7͍��|��W&":�ݚ�Н����F��O��;b�-�2��;�P�t�5$f��_Ub���uQL+��φ��<�6����:��1=���N�KRoY����#�`18vP�� ���Jx�y�Zgl�fb�l����t�h��W+��W��Ɔ �������4�Ք�R'cf���³5����U��+�Xa�H(�˕�Eo(d�J��:�����nސ�ѽv1a{J�k�Vx3G�������S�CП�HN��R��?�d���&�N��	�Ȓ����vm��.�g3Zdj�t��a"�6�m��C������06S��^����$����2�"�1	�<����ߙq�|�����Z��㽕���䕠�s�����혅vº�w�⽒���M���o�G�m�?$��̼�K���Z��㽕���䕽v1a{J�k�Vx3G�(���27:��`.��5��C�)���t�Z����S�CП�R��X鷴QW�w��fD�Ɔ ������&e��c���L}���1LdO�{PH�b_�C���#<x=aUh��������-VL��y���[��,_���p���,@��a��NYs�����4$�[�l��~��R��ƿ;W ��.���:�Nz�]'\gWg��	�Z�kfc�_	�Ƽ���8|bs��2[�a��o���H�RtV�^�d�@���GE�g�������(ӈ���m�r����*qA����6\�4�@�� �-j�1tSjv��
�t��T&���LQ�/81tSjv��H�����4br������Ľ����Չxv��Օ��qvdЧ^{�j����'�����Z>ؼ��XyH�RtV�^�G:w�䖬n���~�����q�ZLN�	��MdGN���!�`�(i36�ZV	�	ҙ���˦G��d�@���G6 y2��R�՝� s�#���k$ �>=���#䖬n��؂�nF���<�W�.�P�	��
�Q�}���%>�rGO�D mWN���%>�rGO�D mWNHN��R��bP�63Z�t�5ߧE4��Fr��j �_�ȇL�X Hz��0�Jw��3�+=�4o���+��+}�K=���e���Օ��qvdЧ^{�jM|�"D5�O�%E#P��=m緒1d�;q3�)�U��)���Y;e�iK!���d.O.C��|#HK��A(�c���_G��Hb� h�ҩΟ/��mS%y�W�CbE�{_8�Y��=�}�Vݨ��}Dq�f�	�)��&ghRV��R���P�|T����{7�H����8���O�υ���YN
��)e#j�o����:5A��p*qA����6\�4�@�� �-j�1tSjv��H�����Yu�������&G!�`�(i3�I��� g�����Օ��qvdЧ^{�jMdGN���!�`�(i3%Q�[�J����˦G��4br��6 y2��R�՝� s�#���k$ �B�'��a����aGl���nF���<�W�.�P�	��
�Q�}���%>�rGO�D mWN!�`�(i3]���-_!Q���ŴIh�5,Wlr�r%)cA/�r�]/2�ݚ�Н��ߎ ��E�VTҝD!u���o���F������}Dq�f��	��x��ݚ�Н��ߎ ��E�VTҝD!u��nF���<�W�.�P�	��
�Q�}���%>�rGO�D mWN���%>�rGO�D mWNHN��R��bP�63Z�t��ܐ�}�k��{`.~��No�ߏ��T�4(���;��|BJ�U�� �X�G[�wE�=p���4br����3v�qh�5,Wlr�r%)cAQ17�b�����d���!i�/��mS%rƂ�o��+h� ��6j�"HsP�����X�G[�OL��qt�Z���#���2=��h��IX0F�MV�ҁGG%4vkz���յ[+8��r$ɓǃl[�Ƶ�1tSjv�>F��3��mlr�{��|e��0�U+�qbp@��߆�p�h��d��JXl'�T��~��Uг�|<;�jmT�#�,l����M?��y�!�`�(i3�}�P6@��e��>��Օ��qvdЧ^{�j@��C2K�ǽ$�!b����#�GWW�<om���濫�L��� h�ҩ��H�������M��2��22= ��v�8:?�'����-����!�`�(i3}�1�Hz8�ZF�*�Gx�����}Dq�f��	��x��ݚ�Н� ��4E|���Bf����{_8�Y��=�}�Vݨ��}Dq�f�HN��R��bP�63Z�tHN��R��bP�63Z�t��Ě����E�i�m}6O�D mWN��ܐ�}Ĉ7NU�.j��u�Nb�BHn̐2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc��TZ��}�S*�"�=3�Ҥ�P�X��������3R��kѶ���� ��&��h�?i�H��}��?<����G&�;���� ����}p閭3u��N�,?��΃���]�X�ֻla�oZx�i�xx�j�甯�[���pФq�Ǒ)''��m�9X��W��� �_%B71Ձ"�Ĭt�'�ǅ@s�-6��P�%Ae!�`�(i3<�6�Q=������Kd���{J��&�)HVi�pz��AY���Z�@���v��d�-td'�I1L�S���%�4/�p_�g�P���V�Wb<�..�4���ho7L��2�"�G�p�Pڹ��/^�w?�d���&�N-Y&yo�q��=m緒X�X�pF�{_8�Y��=�}�Vݨ�ʥ��F��|����"�`Ec'�\Y-φ��<�6�@a� ��fFMqlgd�G}%����3f���K��M�ZP�����V��)�)��H����Qw�c4~Nr_�mS8<�n�ݚ�Н�ʬw�S���q9+t�}�;b�-�2�k+Q�h'�Ȝx�5W ��̫(� h�ҩζ
�t��T&���LQ�/81tSjv������$ɔ9Q<ϯXr&ߜ����>05H~
�:qEp�;�P�t�5fĉ>99��A0ok�׹�x+��IhШ��+���Al+�H�A[�á��'G�+p�Dʾ��6�o8:4�I���c�90B3v�A��{y����i�q,?5q�+�#4��F��8M�H����Qw�c4~Nr_�mS8<�n�ݚ�Н�2VP��Ѣ2����L��my$�N��o�/���;�Ra])n#���^a�nu4Bޗ��jw�	���ݚ�Н�y�}�6f&r#o�]�ʄ�<�i�������M;C��!��iKk�������J*�Rs�08�b(����<��#�!�`�(i3�j���%�|�;�ƇT��J��sr�l�ԝy'�fĉ>99��A0ok��$f��_Ub��7��G_��$�)�vx'X���5����'G�+p�9���?�(�JZ�Vk�;��|B��loXBȱg�S>X;Z�˯��R����e���Wƍ ٻ�l���M���R��ӟ-���4�&����Z����`	p�=�3Yj>�B�R���$]'\gWg��	�Z�kfc&�2���� ��b�FP&�r�@|�TԼ�\�v��_�R�GO.C�U��B��-����A�;�����\�5ｵ����;�jmT�#bs��2[�a��o���H�RtV�^*�9��.����N�eM�#��}Dq�f���NƥNoz��KUq՝� s�#0�ʂ�j�Ï��	�l�lM�3 H�RtV�^܌;���'����u��r���'��o�u:��_x���O����]�!��	Ǹ�y85��8��,	iL�*dgN;ۍ����$9���Z��o�^��D���:5A��p��(1l�jG���Z��o�h�G KH�F;p�	%Ɏ�Bi!�`�(i3�ݚ�Н�-��)'���N�R���Va�irl�
@\�h�5,Wlr�r%)cA/�r�]/2�ݚ�Н���������ۥ�Y�m���NM���!�`�(i3-6���[��<�p��Ar�8w�B
�:qEp�gdq�_x����Yzw��(4G��>��e��>��Օ��qvdЧ^{�jMdGN���!�`�(i3>�Q�c6���*(H=�ƍ2���l�!�`�(i35���u�L����˟y!�`�(i31���~!�`�(i3ʬw�S��ht��p���j��8�u��ݚ�Н�$f��_Ub�F�S�1 �$f��_Ub�F�S�1 ����F��O�}�	76�&�φ��<�6��}�6�nq�Z�@���v�_{ޣ��$7������φ��<�6�@a� ��fFMqlgd�G}%����3f闶P���`�3ޕ �|#HK��A(�c���_G��Hb� h�ҩ�EOJ�uxm�7d��2�4.K7͍��|��W&":�;b�-�2�k+Q�h'�Ȝx�5W ��̫(� h�ҩζ
�t��T&���LQ�/8�@�����2
xH��!�`�(i3CT�MZ�\�XƤ5_��,\���*s-�e�2>J*�Rs�08�b(����T�\yb�����Z>��A�$�|��'T���+�L�F.0D�	�I���_
�u�����|�G�p�P�C������H8Џ�Ӿ���yi�1tSjv��wӨj]h��J��sr�lv{��lw	!ݞX�����}Dq�f���Ě�����}Dq�f��5ߧE4��HN��R���IX0F�Mn5�b	���J��sr�laT��3G?�d���&����*�����E��h���O�Zj�������1φ��<�6�@a� ��fFMqlg{y����i�q,?5q���D5P��wFlE� ��'ž1�|�'����u��r��i��H�p��ic)�̩ƍ2���l�*�9��.�ԫ�&Np;qƍ2���l�����g�Z��3��a���!@�f")u��r��܌;���'����u��r���=�$���Ly���Cʬw�S��ڏ"/��z�>�Q�c6��?��!�6ʬw�S����}Dq�f��5ߧE4��HN��R���ء�I��߸��S�Ȍ���D5P�����+C�!-T��T�^���h�.k�mb�&��ƭ������xO��̋{b62�tstF�!��cܤ|�)՜�45�[՚1Dq��P�<
[�л���7Cw�Hm�̶^�+3���e]�#�?4�s_o#�{�U��)���Y;e�iK!���d.�% ��\:Fa�7�����~�L�D����C#/<���q�r$ɓǃl[�Ƶ�1tSjv�����,<��c�!{p85E�g�������(ӈ���m�r��������x���^a�nu4Bޗ��jw�	��C#/<���q�
�t��T&���LQ�/81tSjv�k��u������}�Fe��1�:��g�XW-#��=���;�P�t�5:Ha��VK�;�P�t�5E�xa�/ݺφ��<�6�2VP��Ѣ� (<ݐ�k-|���vG����и;2z��
�@h�5,Wlr�r%)cA��z>9�R��d���!i�%ؙ,{F�}�1U��VP��t�i?�i2�.[W�w��fD|�O�E/�Ĳ�=�Z���^��[�n�2o� #�����M<E��'Z*)�?�R��n��h
:h����t�h��W+��W���ŊPTWo9���gѸ-���֫IX0F�MV�ҁGG`5:�����+�^n=\f�5>����Db^<�..�4��<qs���|#HK��A(�c���_G��Hb� h�ҩκ%ؙ,{F��#QSU:�����|e"�O)�b�c�!{p85E�g�������(ӈ���m�r����̢k���F�KD�Vr[/}>5��0�B� �b�Ъ���l��=�O�-v�*_�mS8<�n�ݚ�Н��%ؙ,{F���\D�E��hW��ڬ!�,���6+�<�6�Q=5����.������w�h�8Vb5����%>�rGO�D mWNHN��R��bP�63Z�t��ܐ�}ī��K��M�ZP�����Fz��Ԥ���엝�����L}�]���4x;΂��m9Ϲ@��2��w���.�
���t�T��?E-h��`f���sC>��Ӛ��S�J\7�p���"Z�v��!;�jmT�#bs��2[�a��o���H�RtV�^��~Щ�%��v��՝� s�#0�ʂ�j�Ï��	�l�lM�3 H�RtV�^܌;���d��-��!�Bt�wz3��0��I8�ѐv2�_Y�d��o��b�Bϱ��z�
����{�g=_[�7����닓.�`�39����6��ݚ�Н��L&�Ǟ��W�VL��׬��P�|T���nT����
y���^��D��G��q"Y��;����rx�pj�d!�`�(i3��Q7lY��u�M�Һ����1)uם�!�`�(i3�5ߧE4�퉅�%>�rGO�D mWN�Fr��j0C.�>��VaT��3G?�d���&�<��vQ�zi��Hy�GE��R���H"X�0��n���l�IX0F�MV�ҁGG%4vkz����`���φ��<�6�Q١Ӿ�$	��1�h\���F�`yx�>�+X�M?��y�Bz�;{/�>��]#�y�W�CbE�{_8�Y��=�}�Vݨ��}Dq�f�Y�)�}��EXs70��nF���<�W�.�P�	��
�Q�}����g�Z��3��a���!@�f")u��r��܌;���'����u��r��a�F�������Y���D��3��b�]결���:$�O���jF�ཕu�_�mS8<�n�ݚ�Н� �#0xg�`�I��Wz}�ἱc��-).^QQ�b��~$�
�:qEp�;�P�t�5����l��~��?�kv��.V��:��������kB�����X!o%�ſ����O?����<�5�>�?�R��n�K��$�<ۧ�: ��ao.\C�kFGˤ]u���:����
�ݚ�Н��>���Dl����|�b�и|��?���a{�w�!]��̍��}Dq�f������!�`�(i3oj�+p�K�J�iN�SE�g�������(ӈ���m�r����fĉ>99��A0ok��$f��_Ub��7��G_���;�P�t�5�׹�Ӫ��*$���A����ƃ�Y���D��3��b��-��|^a�����Q١Ӿ�$�XƤ5_��,\���1�Hs�k���*��'���9���T�Q١Ӿ�$w���	�e���0��Qܓ'{w#/ B!�`�(i3!�`�(i3$ʩ�})��W��CX-+;X���X��ͷ(�-��]a;����D厺��+�XƤ5_��,\���q���7?�R��nI4�p� ^�b��v݋N�����AS�$�[���G��f#��O?���#j�o������6Bj�!�`�(i3!�`�(i3�����z!J��/٣��q8h��^�Q[M��P��#��s�'	�?��[��羹�He�-�c��R:k�ڛ���Ο]_Z鎬�����	�7 �#�E ���� ��M�#зq8�Ј'���Xw�P���w��a�e56<�5{ΖM+����+�J���q���U��D�U�2Y��i�p��+�FJ�9��V��Q]� _ό���.�@?d�s�8KFmғO�4}`L����D:�n`5�fK�\w��0]\o�LCd�|�w��DK����$���7s�9���o>��l%i�-}�
�?�v�-���w:���z�Ji��d�٣��c�A�L'Qī�*pY�M�l��S�J*�Rs�08�b(������l__��E� )�&��"X��[��Q[R�7�$��Xo��� ���Lk�Bgt�#P4];ˍH��M��=�&&ĕ^$&�	�s�{܇����O�յ[+8�a�)��Ƃ~6T���Q�x1�~g_�,\ަ�It��+g[�Zt%��m&<>��%��JU�a�(�n����62�tϛA^��'T���+M�Mb�:u�w�vG�q�:�&����#|�1�0j��*������Э~���V��2
L.�X;p`��3
�v�v-}�	mp,��_А#�<om���'$W$�X�t����}�(�
4��c��^�
E����d���m l�o�&�C�/w�x�P���E�`JcU!�`�(i3XO����0¤լq��/,���9^-��X�0���X�q!�`�(i3���)�>�)x�?{���x.�Knq���;W��ZLN�	��f�?ǉ�=@�#=���ix���!�`�(i3��ԫrI�C�i�4��v�(��.��dLG���6!�`�(i3���K�7��1۳ఋ�ݚ�Н���*dy�ZB\w��B���!�`�(i3�)ύ^��R�^Ƒ��f�?ǉ�=s���eZ�c]��E���!�`�(i3Q)��Zl�z��SR:g()��ikp���H������7Pr��ġ��,�a��OY�P�CQ��Bރ;�{��C�{����K�7��C4%̈́�(�y�|����x��~iM5/�S3 <�X;p`�M���ʄ?�k�V�?egE�@��i!�`�(i3-��,%>ʴ����қDO,\ͨ܉p����O,8�ݚ�Н�7�N�-��#l'U:�g[q�vG+|�<竷b��"&�_~�:N�4�0 L?�p���@Z,�ttT��Q�#<4^�>N0Θ��ݚ�Н��0V32;5�-�����4)cq�vG+|�<?V��j�cc����L�{��%ў׫>V��2GɎ�#���?\a��4�czZ��������[�D���~�ߗ���@Tvs�!�`�(i3�$�~c/�R��ŭ�.
�:qEp0���Y$���/ӳxW8�8J�|9 �P���R�A��4�h���!U�020�$�~c/�*���J= �P���R�^=^���3!�`�(i37�_M���{�� ��YOZ@��5�h�ʪ%��18�$��`��UB�L5wG�!�`�(i3��2]��ٱ�R:k�ڛԀlY�{:fh�3�w�	�|�s�Õ�M�<���{L,8ԀlY�q-�~_@!�`�(i3�[�H���,޷��u�2�1�9~F�r�t��b���չ�Ad���Ô�b��N�[\�i�]���B��E, �c��ΞOߙYĸ-�4:� �
�	(��7��F�dHw(��ES���v�8:ۛ@W:���#���FӪ�c�g<�j"Xt�F�)��#L����@� ��X�u�%h�K��(�%�z��I��s�*2��3��Wғ��7��&���oC���T8e�i�������ᳮ�T���t�T��?E-h��`f���sC>��Ӛ��S�J\7�p���"Z�v��!;�jmT�#bs��2[�a��o���H�RtV�^��~Щ�%��v��՝� s�#0�ʂ�j�Ï��	�l�lM�3 H�RtV�^�$XR�QܛOcOZail������&G!�`�(i3��Q7lY��u�M�Һ���BO#LB�q#a�_�̞��>��3
�v�v-}�	mp,��_А#�<om�����M��2;!�`�(i3�5ߧE4�퉅�%>�rGO�D mWN�Fr��j�p���"��NwK�"�Q=C&pm" <{>w�\�S�-D�I��L�@��8Q	��+���XƤ5_�J�	�LÆ���#��k���Ϊ�iIn���I_�1����!�`�(i3��7I���aT��3G?�d���&��J�p�k���\�#�k��m6[��!N�'�y�G