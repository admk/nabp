��/  ���B���+QZ��J��S���J��S���J��S���J��S���J��S���J��S������c`�ĶD?=N��J��S������!P7TǱ�J���GRT����<�iQ�����3�7Q���=O ��-K�趹���J6�qQ��J6�qQ��J6�qQ�2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����VcR �z��)��\�4�s�3f]Ǎc��s�lH���G$l$��<�lVщ��~��1�:�Ω��W N��|C��#�N' ���x�t���E�L#uc��WŬ�+�-ޗ(huUP���*+��`�<�R��
�n�T�+F��W��`h��>��ׯ�=>)m��U���T���딣0&_���X0���2|	p��rw@	@us���\���Z�
ۍ���yq�`݊�|���"rG�
���}�\�.�DV	��dU�;�\��^�� ���K�}M^UQ�S��)�e
�9��Ax!P����,��*�b؏�@�~�S�`\��Yi?��n;�|-���g]����g�����fP����IL�+��ץ9�^kh�u��<��T��� �}+~�8Ó B]�pE(���B��|+��@-�-'P�e`b�T=폳�H?o7\F���r��RL�a)�ƞ��U<N	:.���n��{�'����������7C��Hq-/��@�]\���<��9�`J�=�OLl??�L��y�����c��(r���U����D������9��m�!=�y����h�}jh�6g��+��� ���k�o?�M��;]�Qs`k�sǈY���K��j�r��!���<< �sN۪�c�	u�~Rp�,k���%k�&ָ��sE��D�őⴔIꈸV�MT7xB2I�d�HnULkIh��:h
�[ϸ��W�A��S;CM���2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc�# c����2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc2�����Vc(#`��Gcp��}K��f<�,=K�F~�?|�[_X��ˆk�=�r���x�i��p�7��Xi9�
�ѹaB��Q�//?�s�m/C�H*�m��/2�ޅ���?�y��h��ؒ3����]ͧF���y: ���s�JFAa��Bzb;ym��+a��ʁކ�+��T��C�NJ���1�:�Ω�*���g S��/P�p�i/-�#�v-~x��䂁!�o��c��(r���U�ј2��<���ħƿ�9c��?��J��(����5�2���[@%����nEA��"0�qv+d��q�G�+��T��/o��إP�e`b�T=am�������V�2�Ct�z&��ÃlO ܅d^�R@Κ�2���ei����L�IÙ=�HF���m¡;-;*�7��ʐx�?ێ
7�\ZŴ�(??a,����\{F˯�+)�Y-�E�f��Z�>)��p40�zɈT^�`T�W�88�;矷	�gJ�ÃẶ��Ϊ���Jjz�I�~�џ�.���hGD@�F��q���i��I<��fҾ��9��a
�+��8w�=�J�5�o��C!T*Y�{'%s���'����F�r�f�t��6��	���`y������q��ww�=�J�5�o��C!T*Y�{'%s���'����F�r�f�t��6��	���`y����q��G8����<L�|��]���c�A�L'��!�a��5�%]���a(􆿳����^��+��%�k<� -���ݥI��w��,������;�<G��[���ei��"X��[�I�!"lR�^Ƒ����"X��[�d�a�4$�f
�[$��o��C!T*�q���U���d\��N�By3��<Z鎬���������o�	����}��S�)37J*u>����CΊ�?��[�<��z��}�\w��0]�\�LtF��o��C!T*�����2%=dϖ�i�@O�x�7���q�©���$Z�5�8z�E�^^������kK�N��ī��r��X/��4�q�:�"��yȯS���Qߵs<��7�m��+Ȑ E�������?9���Z=%��k3��a�
_g��c���C�x��T��=}�ŕ�F&|S���T�\ ��3��h=T���GZ>.�0b0T��@+���RY��B���M�I@1���t$I+�V�6IWJE�YY���F;�I�e�,��[�9q�Y�{'%s��.|Z���I7��-5��6��	���`y����@����gG̓���#/��p8�(�E;*�}Ւ�~ܔp�l
d
�3�x�. k�|6�8"j���b7|#9���hY����r��4V�H�%ht[����}����g��V)��X�F�r�f�t�8��#��cx�S�����S8�/ #O�)R�^Ƒ����"X��[��Q[R�7��z�h��47�k��9�c_����+�˂߮<ur�<Uee�,�Aٺ�H�'@�"�Q�4V�H�%!.<ή�$���N����]�u�L��ۊr�S�ML�j�|�{');�OA�uW7s�9���o��S8�J�]=��R�^Ƒ����"X��[��Q[R�7d�x� �q�ܯ	�J3���X�/R��rs�i�� ��*b��0��E|�,�CyW�f�tR�wX��}�
�?��V.��(�t%��(��+'���Xw�j�7��ct�:��RE��W��_�ړ8���/����,DpR����Uq4+��]�!��	Ǹ�y85�����څ��;�¬pX��g��U-�e,%�0g���[�=�5x�:�d���G$B�E`^n�&�
_�n�@/%{�;����Q��ǺΕ�f�f3'�g��U-�e,%�0g�������DzL������B�E`^n�&�
_�n�@/%{�;����Q��ǺΕ]I��>��8���/����,D�=P��[:=ȟ�H���
��D&e�2l��4�i�2�X&l����_::���`y���ψ><�'2!2�X 37�˱�5_=���$�4�\_�=@�G���r�ϸ��#|ShI�ˋ���Mei|��sD�hV�\w�4�	H/�"�����ʛ�M>#�!�`�(i3Y%T��BP��&��J�UG�s���#�n�%�y!����-!�`�(i3�a�\����8x<�A!s���Z����Xc����L�{Y%T��BP��&��J��\��;�,S:H��+܆} �S�
â!�`�(i37�ܥ��2�A�Jr���CVF��g�M��p|�\m���X����)�ak�m6���D	��U�l>o��|���bǬ�=����������622��fH��>d]=]A��O�T=�4e=��-Y�VN�=�ԃt����}ꇐ�622��fH��>d]���+�J��U<o^.K�}/��<Ӭ�/�"����J^L���I�PD�naзq8�Ј)w�<�_N`E�cvR+��}Dq�f�(����O��9�JzM�E����F���8�TP��@E�`�8���&��#�@�o0�&�v�x"�,�>E��ʆ�In��tT?�7G|`Y��j3��� Q�N��*lOO_NK8��40=�4e=��-V�׍A���}Dq�f���<E�f��V�mK�b���G(������8�TPO������=��w�[�4�Mei|���)C1Ew\w�4�	H/�"����0�:C&e�!�`�(i3!�`�(i3�a�\����8x<�A!/�"����kU0F�o!�`�(i3!�`�(i3�a�\����8x<�A!s���Z����X�B�r��!�`�(i3�a�\����H�:"�\�(�6k�4d�����͈��}���i!�`�(i37�ܥ��2���kܪ���*�LNm�Zt%��m&<2O!j����x��B5�!�`�(i3x�]�V���M�K�=g�H{g�q��������b�Xϋ?@,�Xʚ@h"�,�>E��4];ˍH��!�,���;���2[����|��1���Wʁ���p�B�E�!�`�(i3���+�J��U<o^.K�}/��<Ӭ�(�6k�4d������z!�
�W@!�`�(i37�ܥ��2�`e7��9��×�>�濖��#�(y��K����!�`�(i3�E����F���8�TPm=_g}b��t�����ܗ�J���� ��A?Љ'�-o��`%��)w�<�_N��M��+?���C&��>k0��w�*�fBg�!�`�(i3���+�J��U<o^.K�}�d	c�b��8���&�Q�$_���]��3a��!�`�(i3=]A��O�T=�4e=��-Y�VN�=��`
 ֢����e���W��]��3a��!�`�(i3x�]�V���t�����[F�a�+�6�5�p����Rܖ���B�r��зq8�Ј)w�<�_N`E�cvR+��}Dq�f�(����O��]��3a��!�`�(i3���D	��U�l>o��|���bǬ�=~�Y���(���8���VZ��W�d�"�,�>E��ʆ�In��tT?�7G|`Y��j3��� Q�N��*lOO_N-�4��j4];ˍH��E�(��<���A�� ,�ttT�r�pΚ�w] n2ϒ��[����r-����8�TPO������=��Z��( ���~*񇦳��Hw�6ٿ����зq8�Ј)w�<�_N�b���VVA�ڦ�c4���ɺ�y��k��)0��=M��LO�|43��52נ޼��X�B��+ H!�`�(i3�E����F���8�TP�}O�6`-�b��Χ�����BQ�.�`��SxEWI�I+�!�`�(i3!�`�(i3"�,�>E��ʆ�In��t�hFyu�.��J��ߟ{�����8n%d��z��BB���#��`'��e�x�]�V���n:�t�c{DJX</��}Dq�f��D��[�
�:�I���G!�`�(i3!�`�(i3=]A��O�T=�4e=��-�ĕ|G���t����}�[V�ct�!�`�(i3!�`�(i3!�`�(i37�ܥ��2�A�Jr�۞��Ѵ���t����}�-O�9�nd_p.���R`!�`�(i3!�`�(i37�ܥ��2�A�Jr�۞��Ѵ���V�52SG���C!�ªj��졼�!�`�(i3!�`�(i3�a�\����H�:"�\��|#HK�����\��w��;�����e��H!�`�(i3���D	��U�l>o��|��@	J�!���}Dq�f�!��I\+��M�a5��|���瀆!�`�(i3=]A��O�T=�4e=��-v����]c�VA�ڦ�c4#B��F�7�ܥ��2���C�0��(����r���� �G�|o#/GD@�F��q+�#�!�	U�E~�˲�<�!�d�<6E[�:x��7JS�����,MLG�j�.(Wx*<�6�Q=�;~����%ho����G���r`
 ֢��FE����墝{l�f|�t�K��0�!�`�(i3!�`�(i3!�`�(i3�;C@����3a�LD�P��Μt��/N�M�O�IQ���}/�"����Ʈ芪�x+�o��C!T*p�VU��J!�`�(i3!�`�(i3!�`�(i3"�,�>E���� &N��nF�d����M^�{�W�Q�
_�J�g�J�LQ��w�mK�#]2� r��w��S�)37J*u���{��}!�`�(i3!�`�(i3!�`�(i3�b��1�K�+��o�.@��A�OH��*Z�h�TD��L���2��}��g��9|P��{l�f|��rs�i���YN���G����exa(􆿳�xE�zH^�7�{_8�Y���˂lq�㜯}Dq�f�F�d�����r<K���J�LQ��wEOJ�uxm� r��w��S�)37J*uc�A�L'�t�O#��XvU(�8���/��}�Ш���my$�N��;� ��b�� л�w-H�.E�^��\=��
i�c�r׽v1a{J�:�r�7��'���Xw�j�7���N�v�1�����7����`y���ȓM�Me����Μt�'�al��p��B�NoSƏw0���8��Q<��z��}�0z�cUL��լ[po�uYG*٦� 7�v�ԯ����fbK7͍��ճ��)�ȓM�Me���섫�So#�'�al��pz��+��ݘ<�6�Q=��f������L�}*2#ԷN�ڿy?"S���0S&",f�e�0�؍�3Ϟ��M�+,[�� л� Ƞ?�T8�� л��d�Q���S�"���=�R���=�u@Ý��},��X:���v�,,�kQ�Ǐ˨�g����K���=
��P��bE˧�<vr/��S�s~�k<����-Ի�弳$��P�!Ўx���-�z%8;����v{:��h���1���N��X�'�f�E�k�8�"�$�����o�u�/z�u #��Mgs�4�H�O��	�� ��Fw"��Aњ��f��>�%Mg�� л�G/1avQ�e�b�����,��Z?m��r�գ���VRj8�@ʚ��X��9�����Ïb�}������c�.D�"]�ϓM���o��C!T*p�VU��Jp��T�����hy�%���[��S�)37J*u�,�JL���*��c�d}];�SS�qL�\�Q���}�+�^@��#	Ͼ7�Z#^L�)�4)	���E}];�SS_�⥳�"_!�`�(i3!�`�(i3�� л��У��a�p�탯;\߰ �Ye�]r��8���F{�grT�i`YS���UP��v��!�`�(i3!�`�(i3<�6�Q=�U�"���M]�B��5.��$�]��tK�"8�f��>�%MgY��j3���d=���ǄҋX����L$�����/���NM����s�٩��8bq�Be��]�!��5��E0�ƺ'���g�{ ,Cѣj�k�-U�P�d���0\��1���FM��`��\n$̱~"��>d�c#�'����1���<��$��tf�E�k�8�"�$�����o�u�/L=x��gO�+�-���qJ�?�̿��{Z�|bQ��� Ǐ˨�g����K���=
��P��bE˧�<vr0�����i�é�I���z�S�*��iMOPԙza��5N�ʡV�l��� л�/�ދ}Ղ�� л��d�Q���S�"���=��
��L����1��in���� zԻ�弳$_N� ���ui�X\�̈́nlH�I<�6�Q=�w�3����f
�@"��g�����R��H�O��	�d[��K�pHj�4�\��ލRC�|�"u�ۼMQNv�2�^��)('���Xw�����C���������C���/S�)37J*u�,�JL���毘3)�:�6�5�p��nz�����:�r�7��'���Xw�����C�������ڥ9��[ʫZN��ҋX����L$�����/�����zQ�.�`��Sy2�H	�?��ҋX������S8���4E�]�V����ft]�c%͠�W7�v�ԯ����fbK7͍��ճ��)�ȓM�Me����Μt����a�kEӮY�E��vNd�)i��Ŷ;���])���/�Z鎬�������(���yf4l!X�t�<�'`ٲ���=������T�\ �͘�f��p�b�z'hۉ)[텡#����Mei|�p��D,L�Y�U��Y���D��L��ȓM�Me���᜶�
2��t��L̿��$|�/|�z}��Hn�[��!'|sI��w��,c�A�L'�t�Otj{%��ߛ�8���/��r�;`��2���<SM0.��~��Ѿ7G#+�Ǘ0z�cUL��լ[po��vf���g��U-�e�dfa���W���n�)Q0N�2߄�%=dϖ�i�B0��O2��p-!]Й���9�{�Jj3ů�/�ۖ��WaU��4��}�<�,3@97��+�o�J:l</�'.�w-�G��HZ��_V�VG�88�;矷��N�����?�d���&����q��w);�OA�uW!�`�(i3!�`�(i3�s���6`� �3�<�G%�MP3$�x�Wt!�`�(i3J�a$�Y F�*3����D�`��p��e;�!�`�(i3�2U��`U��lw�_:3w�⽒���M��ҹf�f3';��|B���r�����M�Q��#�?f�̗���\�rҖ�A$�P�&�2����{y����i�q,?5qM�>Fr����7|)�`����l��!�M��9�a>*<UB3 �~k�%�������&G!�`�(i3�+?B�OA��At��D+���4Y9f2Pih{?��	��٨R��#H+�
�:qEp�;�P�t�5fĉ>99��φ��<�6���(����
W�Q�x�[�g�DPp�$�ҞC���!�`�(i3λF��|�o��_�Rz���n Hd=��¾ȼ!�`�(i3�璓�c�������t �[l;M?��y�!�`�(i32W���R0�����e�����n^-ݖ.�T�w���1��?�Āsf�e�}s�dKa���z%t��#-);�OA�uW�H���~�����l��jZ\C��>CM?��y�!�`�(i3`�~Ӿ�1��?�Āsf�e�}s���xᰪ�!�`�(i3Z��H�H��Bϐp��!�`�(i33��0�����m�#Y�N��b��?�+�ϸ�i�z���v";��H7�: !�`�(i3�5ߧE4��!�`�(i3�5ߧE4�퉅�%>�rG߸��S�Ȍ��8�8!s���}Dq�f�ϟ��7�4��e���]8\빜�&� yE֩�sJ�|���F}�	76�&�;��|B9x�a�����%.y�_�V��	��y��2����8��`+S6E���7-K����}�)��E�d�-���geW���w>��Y��d���!i�a��=�����K��ӌ�lw�_:3w�⽒���M��ҹf�f3';��|B���i��ID����k&��At�����~��]z=2�4^��a��ƴDD�����S�@�
37�˱�5�ݚ�Н��,\ަ�It��+g[�\�
�=ĭ,�*y��<D9��\ǻ�g�<��N�Lf�?ǉ�= I���¬B쪺.C�+�ya0�t�"hzf�?ǉ�=��8����x�&��'�ɹ��I�N���B
��!�`�(i3�?�Y0�
˒KtNp����$y̮�K��v ��>b�eIG��Q�q>xױ�u�i+>O���Q��K�&�C�/��x��&^&Y�o�wd��u~xgA���������6%�a¥�������ķ�X&|a�#�I7��-5��5Z��N����p$Z�"���X;p`�;-;*�7��3z%�u�܆�D:����ЊQvN�G-��A�sxW�O٣����ʄRN�]�5'�ݚ�Н����ȍry��	�MQNv�2	P���i�m�T��!�`�(i3�'�al��pGJ�4۶2�\+/��`C!�`�(i3�v1a{J��w��!+��^���X�B�'��a�U�xn�Oq>N0Θ��ݚ�Н����K�Ȃ��苇��Fe#OOJd֯Y��j3���������g�Hn7�(�!�`�(i3B)vظ�u�a�/!O�f�?ǉ�=EOJ�uxm�)7*{��C�ϟ��7�4��e���JS��Ls�G�E
b�+|�&8�,�pב�B��h޻_JS��Ls�q�ށ �~�g#n]E��A��=5���ǖ�!}�	76�&�;��|B;<T�R18��Ժ��F�w�R���y_Nr`e���4)����%���l�v�\�b�;;�O�{�&l����>M_���ow_;O
�ÿ^�� �O��x��=;Y�ۺ�Ub�!�V��u�ct�:��REs�N
�u�}�T�\ ��;��|B���r����+�uB;y�XNAA���v{��lw	+z��D�H�}�	76�&�;��|B�T'[/Ʊ�&UX�{6j�"Hs|��^�p!\ZeY��3Ah	)ޟo�9f1Eԫ_���358�*��I���;E�@R������ix�ag\�'�al��p�M>�I�dBz�Gb��P�����5?�SLq�N����� v��ʅ�b�O4� ��e���]�!��	Ǹ�y85��3}�@�7 K	����n��H���q�	�<�}��{l�f|�ό���.���S;����!��� ��]�!���Y���f,�(����O�:�r�7��'���Xw�j�7�����4��}5ť�7Z�a(􆿳�GAλ�0��Ŷ;���])���/�Z鎬�������(����c�<Q[j�x��]���"X��[�����Oj�i�K�A��o��C!T*�q���U�����h�W;0ǽi�*��]�!��	Ǹ�y85��3}�@�7 K	����n���Øf�oA؈�'�FT��,{��F�"*�-��2.[]ɭ[�9�:��9Kmv�r��Rϻt<� ).�x6��l���:��9Km?s�_{X4t<� ).�x6��l���:��9Kms��hvo���$y̮��Qr����a�+�wVi�W�W��<��W{0`�����r5�8�4զ"5���q�؅��FJ��/��<Ӭ�,���<C��Bn�W���ɹ��I�"&`�A
!�`�(i3
�Rh	HO��-�L��m+)q����h��@:S
�Rh	HO��@hG��gDiYPc�U6Y̲7kICӱ9E����4���N���m��;���g���70��4)�{6�U���ix�ag\��,}	f��ņ�}h$�q�BZS[]�s�%KjB�'�3=�D�9[8{�n�_ }�(C#ƀ��=���a��bǬ�=�M��yr�v{�h<��T�Ѓ�FĠ"\R؅��FJ���d	c�b��R�s���->��d��vVx�]�V��v��K.Ū(T��������Ӯ0|�s����Mр��=���a\/��cg=�èk�n���y�	s�%�.o�rG��XP���X^�ÎC���l���tL:�C�RH�YGD@�F��qW��Ґ�Yj:{b6��P'��?E/6�+��c�4];ˍH���@E�`17T1������Ka�Ġ"\R؅��FJ���d	c�b��PK�k�V�t(]�XnS��z��@���sA�U� ���_V�׍A�M�ſ�lfR	�_�]_�9M��}�(C#ƀ��=���a�`��	4V��_�$2���w��-��3O�v�ɢ������=���a�`��	4V��_�$2���w��-��3O�}�(C#ƀ��=���a�`��	4@F��[�YR	��.-_��hbV�֎c�TL����U� ���_j0��.@.�����gj�a`�����)J؅��FJ��o�C���j)�3H�,�L�RI�miϢΜ��A.e�@H��F��5������'!�`�(i3!�`�(i37�ܥ��2�`���{�L���i���k��u��0�Ej���lM��2�!�`�(i3!�`�(i3�E����F�'n�^0om�i�K�~sȸ�"rR�ԌY&�xL���b�o!�`�(i3!�`�(i3 ���3�ҺIÙ=�H���mL�0ޥ0D���>M�J<0L}�U��!�`�(i3!�`�(i3l0��F��j �i7�sp>KW℀4�H�� ���+-�K�تG1mv��6��!�`�(i3!�`�(i3x�]�V���M�K�=g�H{g�q����Fz�Z�UL3R�b�jT�.��Ad2`,T�N�M5�ˉ�<�F^^g�)w�<�_N�eب�-�h��C�U�cʝB׹[vk��u��:��+���f�.`�G����4�t!�`�(i3�E����F�'n�^0oT�X�ܣ�sȸ�"rR�%��ZJTD�x��]�!�`�(i3!�`�(i3 ���3�ҺIÙ=�H�����*m��kÉm*�-�b�+�